��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c��5�h�:�**$�'�r!�%N7����Av��mrwR��R�<���GjC4 u�E窱K$�g=�d|E�He�<[,Dؑ0�KyO�u�X�Jq�Z}�	�%A�F"�+�Y��
�)j�:���f^f�|�,�B�ϱ
�����bĻ#G���SHҚ2[+���}��~_`�~��]�U�̶�n�p�Q� Y�����#��Y���һ/������k'q��R��@t@���p��Ɔ$�D��2�e����ըeKx��;�)N�F���>�ޗ�l�邍���X+rK�(�d�#�WD��1�G8A���W �+>{K�?��Ѫq��.j�<�FB� Y��+וj
t	���o�/	2R�I�? ���ִ�j�롪\��j�?n02��G�|�����C�������6h��e����ڠ`��*7��������k�/�]�y릚��ܤ�������ַ?f���bשܛ]d�>�-#�W��1��`�(����Z���m�w wE��tw ;����buC�{�P`U�ss�A�8��c��#�r�4�y56d�����J�2��4RΦ�o*��+>%�T2�n��ĉL?�Zj���E��=��]C�oe�kW������E�آz:`��h�I+c�T�
T2�4����U�xݔ_��ih��*���<�� x�PA2�n�-��NP�-:m��-_/$y��	�Ѕ�	��^����:��(W�1ʹ}l���d"$���Ri\�T���7�Y��m#ڮ$Z,]��rb�i��P>{��]����>f�wDTt�=���Ԥ�2K��^d�^pt�L�s	L��X��,4���-av`�kdGb�'��/1��ɔ��)s=1Ͽ�c��-��(m�V���M��)h�����BF8Zm=�%����/*e &���,f�<��Ҷp����%�Z>�޷$W���툛�^ ����,%QV؇7"��P�E��1ƴtge��9�'����!^�eｿ��e>{@��5�=
S����,^�{O�
��]��-y����qFd�<a�u/<�(����5-��,�	s�>`�O$�u!��(2����M]s���C�9�u�� �<�&�����Y�)^WKp\S���,Y�#H����Aȡ m�V�ϑ`	\LP����^����M:�_c*R����c(�M,�M?�w�M��9vk�Ȟ#��\��P�d��mv^��Z���`�nxf3H8��b0�c��8�AZZI��U(mT�"��a�B��h����1��*�'g��B�ؒ���[ب*��qȞ���<3��Ũp��F��|
��o6����@ס*��+,����*)��)���r�BK�D�������;��,�0wG(�261���5-J��^�⫗��U�8�D��|��]�۰8�/�zg��q�����R�K���Y;��]�W�ij�=�A��,s���UZȷ���fM:
~hxjB)�H>�M�c��N����7�z{��vOAV�]���T��@�K�E>7����I��6���;�(�"���Cǭ��90I�d�9α�4���a�3�C�e��l�:up�%�`��Њ�v�s2�ot6΃P3V��Нhdww�F  ���ϧ�����4u�<~�2�T*)\��a����s(.3�\V�B'�ا��lʻH ��G}�/7�_����6��������Q�%�5�� ���&��+Sd��7%��Z��G|����1xj�h�-zu� F%�E]ЪO"�)P�N�m&�Y'��q�~�1^����sw�QF��<Ӱح[�,X(��%�;zF.j`�cm�	ƋV��
�w�f�=җo�D��b��34����_�/9��.�G����j�+8|;�6fT4��[QRƜ�3�k̗s��E�r��]b��=��wIv�E
����Q�w*�aNU.M�4��7p�t���;P?2��s x��q��w֜��ͷ���P�(�r�M@^��ΐX2W~̈ww2�&m�
�y}�w�"	��D� ,�`H�nhx���Lnܓ'�̠�{�����;�%�^	�̯�u4:P�y��	��N�0`Lc߄�Q��c��e<�|K��4v�B��|ٯ����PI���+��V���%��z��Dv��F�����w�������a3���PlI|���Jt��0��e5�KH�f�/)zwa�(w!/i�'D�w�=m�x�F���s�"��'i c����T�Ur��ۻ�5��Ua^q�i3�ew4��]N��L�j���cG[�9 �O��܀�\��Xx�������I��v�&�_^��0�U��F"�ح���K����a��;X>���N
�M�P���G\��D/��������_�5��Q�=!��a��G:��(���4��AAN���N��߽�}�5��o!��z�/*��z
&Pz���8�~�\XZ�O��JNq��8�|�A��@>���~�i_5���[#5����� �������aA)6� uקe���h-
�s{�0 �q�+M�5�N1��]�c)�ۛ�(��ϑ@����	��
^!� N�k%~$Ԓ���r�d��`�$H��l��C�񃉺�o%�^��_��#sd�v9�H%��*�ǳ��L�,�t��E��*�ʙ_Ԧ�&>��j��V�,R�4Ɖo*��C�Nf�4n�Ӡ�K��OmcAq��||�0�'@��"�'"������7�J��ңIz���7�T6�{���$rW!T�uK���a����Ī�畂�L�Q��S�S9C�ۗ�ս��/���$f ��־d�>��n���c��Pu꿻Ƌ��7o��������l���N��Ǟ�N�cT�%>+X�^��U v��듊c/��1y}����Z��_ָ�1'}e�(�꟩Y�>�|��q�P��үG=��_���y�{'(��J�Vr�/��o��dX��ɗ�<tyb�۬����`�!V>���fq����f�/�H�+Rn�����}��gv��.M�x<����,�?v\��x��6���p�N�_:�չ��%4G��2�)n�*��2�ɌHrչ/�hE����XZ��޵�1�C���m��*Q��jt
rțyծ��+.2����P,e���v|){"	�^$��T:��=v��Y���Y�pA�ܞ�B���I�9m+rr��~�[0������?/N��~�R�<�H��W��A4#�Nd����2[�y�{�	�,i$�|)��s��՗�M��DB��
Nػ'��dP���d�̧���V�Gg���+�I�i>1��� �e3��?��\i��D/�M1V�{D=�����^w�q�@�������Y�^Ð��1�q!0�/�6�`	�@O�#w�^���96�݈�c�hI�཮�F��Ma ht���Y"�6�l��[�l����c�Ɔ�O�����hhZ��_�/
�ZB#�c�E1l�_�$��=:{$j�|��T I{ '}��Ɉ2�U�ED=�p���Lb������n4F{	�����^�� r�BG�$�i��ˤ�^]�}��POat#� ^�uWpk���kxp�v�-��wgov&�hfP�#6s�@�-l��$S�s��ς|:=�VN�hq��;h��V�l�MO�t9��K{����I큔8��~�,�J֖W�g'�z�֓��c@±4l!"lN^0|=�"3�=&��,��8'�V]���#������H�f��0��	!F���g`�O��
Y;�Ȍ쁏��|n\8e�b�.Y��?8�LV_���>�����S0!)Z��s������}+}9e [H��n��	W���`�@E��Ո���&�n<���	X14�	1�&��ٗ��,~;��ʡAY��Y�ч �����������Õ�G=�ܮ.Bmd�$K�HId���'�]�3�+��}���V$�G̷
},�Z��c=���?ڝ/�LodcǣX,��e��`��.|����0��t���ԋ����,�t�D��~�����od:�j=�+�B.S��h��P�3e����VEn4��D�vI��C�@t��C�����j ��(�/������Ԅ��*��}��g�����D�L2���U�C��^����#��Z٘��·N�G�x��W�ަ�mY�L1����[q�D�4�`��;��RhGg��!nH�8s��}�T-mˇ4�n�f�QE��!���R�����v�W~���BO*��|�r	�x'm�o6�a��$�h���X2o��}���|�Ej�v����1��n�l5TO��������_���`]J൜?>0n�ӵO�y�� Mؖ��H�~7;^�i;I�G��K��L���2��;Be�x����{���Z:�>�-,ov�����U,�]���Oˆz�48nD�7X�*��H3c�(i�!ӛ��$���W�R���	P�ħ��PY_�[y��Pf�ޤ�:N�j�|���|�@k�]�R{��挓�@��?FI��W���V��঳�4�U2h��;B�-�۞���>�˫��z99��A�뾶�/ЕC��һ�ޤ���,�(Qf�$W��/�9Y��x��A�W[P�RҎD�]�Y�fT��#�9WPyG%�r�'���5j!�SY�c4S퉑S� �q�u�'h2\ǧ��F���;z�!TM̦}t��{�?]>?XAM�%��$3���o��/����]"�C�m[1�3�s�o��Xޮ�:9�Kȅ�uY�StC���%S=�$�ܡ�x$0���c�=�~W�Qc������bD�PN��HT���1֫�F	!��Ă���Jiy�w�E�M�
���C���� ��Yc���s�P�tJ�BBhl;�UBm��3ڔC�����||ԓ�E�rU�H��&ͧ�i��a�Ϯ������[���U�O�_f2D'5�r 𵧰��m�Ee��]�CD���l�S��r��ɟ2l�ޏ!~e�"��y������UI���<�\�W���ﷷ��=�k���;S��K�]A2����uE؇٭���S��t(!���e�&k-TJ=E|�̓0H��UΌ������9�g��_0�E�f�G �4+h#���	>��<�]�=�$���ۼ!�IL� W�e�h��%�v����W�Erp�����OMg?�CC{�~a��,*[���m���cߋg\S���q�bqm_�n�4�����>{�R��+�_^}�3�>�/��j#��t�4D���UVyy��8����{�3ҝ�.�.Rhe���Ѳ�o�+R��تg��.xs�mo��j�K���zG�<k��X���B��_#h�bz��3B�����H'>ͣj���ɂ�R�0�/�uZ >-GO�f������d���sM��d���|Yjt�³��\O{������[�Pw�K<@�.';�������X�;v�����S4Ĺ�������51��Sc��|�0&7��US�0;7�y�琶j�NC�O�iF�8�͌_M����� ,�8%]UF�J�����(�2��=)�+����c,\]�'^��q�i@n���N���`��R�Q�Ҟ�g������gb�����-����+����ꢏx���ô5H���Eœ��
-,�ϗ��KH��"=
4ΐИf�|_�9�W�t;��[�M�����f�w�JI����z/�,xV4��nk��\��!I;s&�M@=��r����n���ҁϪ�M�f�w�"v(��
kX�K��\��t�?2"c��"�Ui�wOZ:Bo���Y��f���ysp���m�EX��2�A�Ui�b���ZEG��U}T,���|{a���<^��lR�d��d&]KM[#�C�D�Z� �K5�ԏ��u�&��Z����cb�ԺZm�C`��X�c���w�6�VMa���3׏4���;�T[�ֽ.���2�]���E�^����"Pm� j!DL'��R{SԼMqǠ�:T}P���0���3U�t}�p/�0�)x�,tX���ů_m�X�>=��9�����`��g��p(Cln [UQ�.b���;��a~F6{إ[i��&�T%N苩|�)�#rF�$f |����.��
~�9O[ܓ�&�/�ڸ���!��~�{a�J�ʹ&Y<A��p��~����f��h<,��,3��>�6�K�-����I��#X�'�z�o7���3?y���� ��i-!�q��9v�Zh�y�����]r�+Wo���������Rꕖ����R��_o��۵YU�	���*zPNև�.S&Äy��Z:��A�_ ���3�Z�Ւ��dİ�C����nr90�1tɦw�VTʓLsʕ��E��*��z�H"ѷ�q|׃G\�}��h�0K��[��/�grRf�d���1�}V�C=��F�yH���6����1��<u���O�Q%��*�V�̏G�#�E�d�$���t^LzK�IV3���L8���_=�������zr�R���y^�ɝD>�����I=�:HZ@Z���3�u˹s��']�؞�W��Q�	�H�:���[!�C�Ԏ������F�,�Ad�� �d��m=r�jؔ��gn^�^H��j}��ެ�Oj����ma�릯)Y�wh�j�o������d�=�����DU�^:���Q��Zc�s���ݓ>��:jn�*|�h��$s���C� x�rR
IHVgE����cd��̍aBYn/kc~�b6�.�,��:�9�8ޜBMgLz��F�����<�\f�u�`9=w��j*3����_h�g]7!rŕ1Su_��:&��<�<c�ȱ��P�HũS]Lגּ81Ƨy�C1g�ݦ�H��zh��"w�u��~@v������p"�t��OK�A��?�G&�����%i*�b=C4`��<�R�E��?<���l��X�p�K�Ӌ��Ln0�h����{wnC�Ǉ�J���/��3̓e�R���K�/.Ơy
h;��k�8�)�H������Z�Y��1�R"{$�`e�q�Ί�S�=}N�cE���/��\�ݬ�&��}���ͥ(��㥧��nM��n��T��O�t�V>�,Ȝ�O2�&��B[qׁ���� E��쨁9%�o_��ݣ�䭧�*E �܆ >�T�k�@Fb��U�-�dNH%�B�;�Y��'5KP�f�r�w�j�t��G�6�z��^��ro��}�ycTeNX�06VQ��(�t�	����8��*]��ʨ��J��Ĵ��_>F��x�sm5kYJG��\P�7X�{[|c䴀��c��F�*�(f�����#@9�zB�h/��R�p���ڈo��Ve�{��M^����(��v+W���M���}I��"śZDi����L��"y���iJ!���-.H� Vpt�%��̝�H�w �����y@�_L�([�م�}���kn퍾��s�y�1�igv?����-!.)&�����.iJ�| �L�ڧ�渒Q� yt�4A����P�]�;���؄3֛vz���n�q�,o7�,�d~Y�խ��mW�y�Qu.�P�
���?~r��Ҍ��p�\�F��S��E�8/sZ�`�Ѕ'��u�U��β���W G���c�Gh���3����t�;c��ɜ��b}��|�K� p����I�2���4���iʰt��x��,��j��t����!c�������7DK�f����w�TuD�T/���_h)� 0L������>Dп�.�D��'"��A�-w��c�KQ�i�D��|�ce��`���ڤ�I����@W��=�^�2�	m�1��mB�w���G�0n����s�� ���#`;����L?"hd��7�fT�O�8L�=�tc����§<P�t�w�\��4�{�"�1�庢@���B�6󦻭�g��YYF�M�g)t�@��DE�Gy'>{��M�9�PE���1/�b�kBq�x��(ꏘ�E3�;��u�'�/A�C;��7��C��3�q)DwO�eV��.�S��]���ST���}���BY��_B���EJ�m�����0��H#��\���ߦ~#�W�Y�|Z��<g�!�W�G�ƹ��������$z���+��f���D�,�T-�@R܆�O��X#+�|~��B�Z���F/���+b/?��[�U���:U� (F��oe/�������<}P5���� G�c������h=��8&�(忟�ur)���.^�s_�&v�H��^G�v���[��T��e7^l�hB��]��(�]ـ�0�y٤��]��� �^���!r^*�S�~`c����J���ž+K�]�O�ޕ�7���2�!�!7-�����<ZR�/S�a�otJ����A;;�MԂ)~����ȿ�]qP�W�9��`8^F�k�4&��-��V��+�7�A��5ֆ̊� �w�i�3��@l��Xa����}p �k�)�u��bRq�Ĭ�����q�=F�gT*�B�܅�T�cH�LB�qҩ�c��[�U�o܍��t�HB�j���P��t���z���I��m'��n��yl���M��2z��҈�.�*��6E���\DH��ઃ���	� ��j�Y,e߸/� .<a�[J���7�"]�#T*+��7ii�]�����I8}�WV�9бR=Ο�E\�)� ���E3
���F6����]Y�nuY��F�%d��N��$T��5b*kSm��ʴ#a�`%NV�@D��J��D>u�J)�c�C^�#E�*�S��Ӵ5�l��)}�1�	?�|��<XS��^^�Tf��+�豚Jp*�W͵�ӱk�8Yg�B��>��K֑$�R�qQ	��,��(
��Aw/]=�+�v�e;�r��T9`�7!l���-!�?(��w|��#ןQ�|�k���ؒ�lJ`��|4�����ӦϬM�/�e퀈+��C#�\�]��=�zw���V�`��L����2''̼��<m�lk��5qBɻ,��G��}M�y07��n$�CپQ10�[��bg��N :��"I
>��3T���H�h��ry�6���B���4�d`�Vq-����ѵ����T��@��6����)�Z���"��<�+�SOZF�-,�R͜�����`�c�雞�I��"|���?&��d���9o�B��Ϟ���ݰZaB�A�HX� ��&�'ζ�^Ҷ�K(���=f��/-F�y=�o��9����W�V�@3�`��̌����M�� !���hJIȑ`��T��w��Qh*UJD��;�V���G��!�wO���1���y���Cp���N�py�AR��	t�O{�,L1��3����rv�/zf��Xs���1"Y��ҡzf"A��v��J9A0�i�e·�c�S�����Wd���I�6�;7�7����a�>���R�D�D���`Q�%x�U��*irǥ����vd_|�9Ž�-�/�Fs.M��0����Ze,�Bُ���|�W-ǎ��KȦsgl�a"�I�I(����Ǯ<�;��K~��I;���UR��
��=ٲ��у�$������s���S:��c�i̯�-�?1Y�T����u������B��H���z2�]�q���_�%|X%�o�>*cy=��� ���	�ɰ�=c�E���#��;��^i�?(�rQjFI�GZ�u�G�<�kί@%�����'D�|�7U���<��j�014��fV����G<� W�$��hDM��ɻ\r���ӫ���%������ޥ�dJh��:8u�4�k,[/0��:R�:�m<�4������\�-�%��A�(�pI"^�Vc߼��M`2�ʥ�n/X�_��p��D�q�O~cT9|���l�.2, )X�����[�.%�������i9V�b���hd��R�ݤ|�a�6 �]>�3��T$�\�f�����(�;�� X��r��y_D����sE�io��a�"� ä|��0�>�[�l�>�aP���{@%�_���]�-���to��T��A� �
@P!�����x4�
��;S��#����D��p��+и2���7㙻Ǽ�o����+�n!D՞��� Ff���D$oyAbc�ݷW�]:I��S�M͓h�_; W��X|>
eAX��Y�������W�o��[@���
����|�i5���!xnN�K
@Xc"9 ��.�H?���;6Y(��@�����ߴ��gˑ�ŧ�;{�&5�����OQ�ڱpW0	B� �5g�M"y*K��Uf+Ht�g�]�� �
����]�ʹ�6�q��t��WM�V?�����g&��C��m�����$
��Y�~D����X��$D��C�K��қ��N�c�.H��Xs<|5wi��0G�$هr&��.w�A�t)(�Dn7Agʩ^�;f��L��w���)�a,�/��՟1qGk���f��d4�z'T�B�R���\�Phzk��V�׽~�U���eJ�ݐ�a�dN�L�&�Q�P�Þt��+S��� |t��H��.�(^ꚉ�$��Z�-C�`:Cb��k�"�n��>XHk���L�X�k�Q���A��^�$sŘ<�����f�:��5�>:�'�:Lz�9���[m�+k�Z��>a���<�k�v�5`��Š.� 2� ��T:{��4j�I�&9z*��A�ꉝ<�Ӗr��Ƴ��]ƙr�^�m�m��5u��M�[B�<�����&���Y:}�6�k/@m��w:��˹"M��=�m�+��]�nY�M	�͕��g�#��}���׀7���l�bJ����/�s__��4ym��2;`���O��I~�/��^���em�dd�"~r+ V�3
mF�+�8F=���r�*�`�4q��%�+�R,i=�u5f�����т
�R�L�Q �5��b�+�,w�(9>C��zŎI�����lI�B]:�Dp����5s���WvL�
p�y�a'�RKGG�^k���U=nI�*R|�l;E�>�����(^�'NP]|���-�)��+�7��NY���(v��~���L.��_�ۼ��r�2��q�<f��ץ��!�+:wł[�_3]�qr�%����a��Pg�r���Ej:@n�dI]�}�5��==P/ϵ^A$���=,�xsm9��b�B|���RS�-o(7�*�/��@?|#J}hf~��������zz� �)��n��n!�=%N��Z	����E�~�eM�a��їDs��u?Iz�#>@4|������,]jП[� /��3e���}��2�H\*��P��r����0T	��1�-��������&S�3}|`�||���Z�v��c�{Ev΀b�{E,��4�<0 /��r$���B	�;~��AO�Lfco\��Q�Qj�&`if�����Q5"�K��"3 �^�J�1}x�u�����{��Y�*�{Fq�K��ks�Jd]�+R( ����$;���t�p�SS�%�8m���7���n�y�Ҥ�z�/��(��ą5�E�*��d+ԩ�X ��7:�0�}O5.��� ������r�2z6mfi���,��)���n^2���vBB���=���Nl&K\i^_��I?�Ӳ,SU�)\�%�J��Y��2�U�䥥����jkwA{YN	����]h�=ޫ�D	�l]��k|oxo�CPXbiI���.��Zk�Vc����c�EM��Z-��#l��V�����n�4`�����*���א+�tr1�>�i�. �Y�O!K�(���F,�4i���Í���_Z�9���(�>?["�щ���v{$xW�0���q0�6t_yq���/i��Ou�o'����XF?�%U0�&��6�.�B�@��)��f�n�{��L_˃����a��k4]�g�5V� �a&�A@��ÄC�z)�N�</��o=Q�[+��TO�i�d6躗a�U��5��D�.8�[[����}�NZX��g6����� ���c\b�qc�k|?��vpb�2�o~�59<t�̩��y��v�ۣC��"T�bo�o�\���5T��M��ٔe��FC�Z�;��1F�sX�WK�%��8p��סf����Y$�����t��ö�#���D���'h����E~k�dm(��0*ʸ4��/���X���6���Ǡ3,���-=$5�P�C�����]����g.�k:�S��	+�I���#��i�iڐ�y�bk��k��T<����3sm�H�o�t� 9�GF��{ �O���hGp�I@V0JhV���Ĕ��9�s�=zO٪=[���y��jcx�N���R��4Z��u⺟��A ϒ�=Kk��}�\ٙ��O�����qC(\šK�o�Ak^���p�/�_���<R(�KR5��f(�ㅉx]�������!�^s�+k��� ���Ӳ�ω�[p^U�� ��
&�Yw����;�e�RE2��@ ǆׯ���x����a�y++����F���i���Q5�3M�4�Z��Y	M?;�g�hy��GĖ��z�$TU��O�vWB���8�Un��ϯ�\���m��t��7�w�z?�l줪\�BzP�+%�K��!��~7��h����L�Q���(��(etYس�}Ve�l���R��|v�� ��QX$x
��f�D̈> �,�����tS	�����(�\wvI�r�`%8b��O��%rGZ�����D�,�I}�d�a��#S��)&���#ȇ��_4�x=���*+�������A��4w���&]�}�y�8,F�/��媟��h�yf�.U65̝$(�^�/)��C7c�e �v�Rh��Q9}p�"]�dm������?Ÿ�;]0�qp�Pn<p�"c��y�,j
,����7��b.C[&��S�{B蝯/x�ԝ��Ȁ^��&_��v�7��.�c��@SL�1�]�A���.��3z��G�����"��4�?/�.5i^<1�S��p���VC)�Z�װ�{��m���d���b���ϳe����<�\ChM�H�$��vP�
C7��.�Ξ�����Q.���e'C�L�	j���a7�r���W���G���]ώ��zS\?��������-�/9�Q��c]h?yH9	n��U�O�_s��3l���Vty��������ŗ�B�&Cʾ��r��5b��1��� ���� �h��,� R�0pN��q%�``a�2�"�w2�⌼L��#�rh�BQ�����Q��5�9v|�X躦���ʎ���c�+d��V���˭�!����=$Ⱥ�ˋo	�i 3�����5d�����7�_�k�ו��N�~���-�'��C�R>�H7�l#��w���M��O��I��pĀ�%�8���ST0�q˃���Z��۴�^��o|T�a0&z��4Tp�7<�b�z�D�f�F�,����)��Ky\3�VM$nTQ:O�bg�g�5��ly�_��-��"�*��QX�1]	r�M(��i��~�E2ɳeI���3=�W����1���}��0�2����bP����pk��!���y�!�ʷV�\��m�5���2�E`�oSg瀲D�g�?
;��4=�],�.6�+{X,[��U�����1�X���\^(��{tD[��׽��V�%PU\՜uP	�v�k���Ҭ�d�������M�N����*�Ţ�*��5�c�=WrS���7Z~�D�����@U��'q�aW8�h��M�mQ.���pR,o�`�p���Ў��Yʹ���D��Mϝ?h-����&pgY
y3Q�pȮZA���q�ւ}�� �F��QN�\(4�M���WyhmZE��ߗ��ޗ����F�	;&��#u,Q�y%��d����A�����iL�'K��J�/L�Ś��ZD>�i#V�'�w��^f*�Cޣ�#zZ�:��~��°~�3f�a�/�S���/����N�{�q�`�5��t
,�#�$+�V!{U� �����|��ȼ�yU����{܋�����>�e8�+��P��#9�����Y3sX��H�n	���9��l���g�l��[p����I����?�S�0�fћ$��6���d�<5LA����+���D]��Sg�Qw�׿T&ZJ�w�^}=���/�O��b�#\W=ep��������۫;f���V�B��E���+�/#:�����"+>�u)0Š(0t�G{k�1�h1���+��L���ԃ�9oD�^�������u�1� �Vj�W�Bs&�?��2�m�^��G��H�hj���N�%����ˑ���M����6�����g��c�:�' _���č�#�t�='�Z��a�Ք�*�G���nn��6�ˀ��M��h� Tl?��jy6>��X��N�:W�d��y[+��-��ָ����x�Q��k�Ĥ�c�n�phJ�T�ȶ8@�ÿ*��L�>��!�^�h���
��$��#�����T�aE������M�5ީx�A,2�z$��'�s�s��������,Z���/�a1���O��Ε��|}N{����׆��+�-�8=�XLj(�pAӫgO�!RtC �c>Ğ�"n��MI�o�w6fZ,^�8{���LU�h�MǨ?Q������}�[�?0�f%.�)��ܖC��|3�:�c[fq��e�r'�i����~��ax��9�Ww[�D̩V�ȭ�q
բk��5���8��;�B
�)��HY׬����a4���]�S|I����;L2�R�:m�f~�c6�,������ц���UZ/�G�u��Â8��������'�¶�gL��e�x?j,<��Y<���X-�7��q�X2f/��x~�\�ii,���M��1�dݴvi�w
 �Q}��r��_�}����\�(H5��]&��������pCA�"�-	�s�jV������(?\B������)U5-e�������!���]�vXt��c�ݴ����j�`%g�#���z��F]/��E�Z���1���;YG$	�ca�22��/t��R�FSh�a�/�?_�y�.'��~S���*�	�`�xF��ߔa�oD�V���~v5G$!�J�:�t�|��{R�hp$�f�N$&����*��H��}�2t�k�fG~2�FB�oV	{��2���p*��Vy��hU1��&� eٷOC�R�t8�w(wkn�ֵ����e��\��i���`0k�o��24���Ա�GqvP^�e��ň�@g	Q&pv��?cB�5�qf�oݩ2����r��	�ȓ��o��G�1b Z�uKҨ�T9Aw�h�V��y�ܻ�~ ���g�(${m�˴N馰�)��S��Q�>��j<�@I�$�`!-{%�\�B-c��FT$s�~q���V�$|yK����+\d�J��
�\cK�I�9�!�ӐX��:Q2��UQ���b��8�DsRVeF��R��)k�_�{A�~���<�Fm�K�d�?�-�|ޜ���Y���k܏Vz���+�w�e��5��L������I��kv�۱@�	��'i�Cc��2Rt�����5R����^|dX��e�ؠ���Il� ��!GM�S�k	��a�̔S+���GMB;����W�N��;��?�=��$��C{�e!��c����Q7~KYuV�=|8]|�����^u1���R'�dKG%SՂ��!�R�;s;�)�����kl����&���\�����i/����\��|����L4�h">	�ő�:j��C����i��T��G��i��n����D��`�0N>�T���K:�1�I,/�G�ْ�:Z��Z��o1��
nQ��@fO���^|eoM[����{�:}H�#D�@���u�Z���6R�5���ŒH�b�m˚Xg[r��g�^�em]���(ā��5��V���N=Q�~�cOS�IU����l�\ ��54+� z��7�8��%X㜬���b����ZM6l�MَO��Sz�^�$y�H3e:�2-/�� q�Ct��%%L-!�x��wk�àJ�vc{\�@�������^�N�6qU� ݍ3JfÙ��)Ǭ(���P=E��4p�U���S3�!���8�{<zq��ޮ9"*��p��8�	vS�?j�u5Bh%r��#T�zFAHt��CU�BN�g��W�[����0H�Uӽ�T}�y^u��,i�<� ���fa�]NG�2~�m��g�r_n� �;�%�]� �
����;H-<m�4	�����.�OЦ���˜���dE��7�Đ��Mm��՘]�]wF��S�ܔ�����;�LQ::����C�xiq��*�z2�@�������V�Cx����2i(�Wt�[��=�.+�<�̊���Ӎ�2���g�d��>_����17:����_�E�E���S9P�A(��r�uV�Z�PO�W�p�_�,�����d� �"�]��v]j)����e�KU��5�~m�I(s��^w�؉���ƿ�U�;�5�V��:��u�iXQ
n�l5��`]T��rg���"P��#���Xf@�V��evϒ;1?��^ G����m�"E]�"���hz	K��9�����Ur_>�����{o��Iu��������s��7=ܯLՓ�o�2���V�������i���K�&<��^�=���Ĩ �oȕ��� �A�F��e*����8�ow,;�Hkg�1�4� �A�Q�&M"���Uz��$�Ό����P�k�m.��g����D�$=��e[G��6�r%	$�]���3jde5�p ����&l8U��s�aD��)j@��g���	��З@s�L6SÂ�[,&~�_��-��M"!�6U��Hw:P�۳98��&���� uĀ�������!P��I�*����T���[M��\����9�~�2Й_H�q��C���l�l���"}}�p�h��hqyto�bj
��_ ��d��ˠ���y!�T bD��^ˏ&ֿ����j�q,|�t�b|O,���1NxAT�QBR>��l&-3j�Ͽq�16�	Vt�pEKF�2- �*���C�eqŁݤN=	a�.%h�7���H�e4a]��ࡄ`��4� qio�ӆyP?�����D��R��K�1%��h�!��-d��e�=^$�	���&[��ٟ{�ُ��� ζ�1-b���Q�q��Lz�IL�!r�����~yנ�d\�{�/����H��h-z�2�w�Z:ǈV�r0�Ψ6���ү��~����W1ʟ�X��V��c��]mf�ʪ��T���� w� �6��RN���h�Q�)�Ha�P?R�*��I�0MmK�U��M����@Q�-RC��_����
@��q9��-P�]'�"��BY�ч����+o漆��,� J$2ֈ*����TS� ����e������ڣϬ��~ܬ�Q��C��*�/P1�d��NɘvՕ��>���� ��
4��SfsZ��C�׆���u��*�Hg�Z�Aw8Ӈ'�XSJ��U�u�k�$��@�z��)B	u-t�7]L+�xV�����E�[�F�;�?��/.r�h� W�d[��8N�B|�����sOa��f�ƅKJ��#1w�߭������u<[-q>6z|U�g�ʀI����_u��p�בs��[��@D�Ч��?;#�^�e TL�����0G֕K
�o��;�h&����9JW���>��5�t9�qY
����3&�ΉQ����y!aS����{3�~�+Ѝ����A-[�2ڤZ;{��<�FTE�1��$�F���n�"*��-����GD�^��s�eZ&�����k�>�H�\?��0�`@ �0h�:���T~;Rt�V�
5���yC�	��]�.�������m����R
����&�A�w�y���%˻�)7�W����	��W�ײ�׻���,��ݷ�T��6��a�3�+�_�n�F �:o�Ĝ;�M\�WB.#�黪�b�<���Wf~����w�4��39���Zs+���"I��V��D�oI"�Z ٕ���RY�e�
g=�n�)k4��r#Ja��1��^)�eh��)0�w�1��s�T��,DD^޳Hު �(���ޱ���܀R��pi}�5�۱׾l�
�D��P�ވ��f@�KaF�v�\�cF�+�|�r��nip�|�9S�3��� d�՞�$\[������>�*��'P���Qs�-ai�""l����� �i��"w
n�`�E~n�r5~�Z���n��A�(�8�I�<g>���yhNA��*�>)!�`Zu�KV�î�	rX)g����]��yf������p{���n�vB��Ss:SL��9#���krZ���:8��%�X!����"f,��NyO
�y�@�	O�Hm�� �i��!�
L�(��I�q�z�"�c��U5c�uC�yO+b-�fz.V�g\��R��/��:I ��F�C�Oe��c�`\����o�\��'��Ni�Ux�4�
z_���S�<[�W{�5��E� 2g��Q��m4D�����H�X�I}3�n���䡧���$S��h�š�Ģ������ԿT��撶X��Pobg��Y�]�p;Q)�:"% ��|R>���"��L"h(S�?�X��,f3�yREO}�c|R������U�j@������~���{��pp�^kBV9p�G�IF�g (c]\�n�w�l�os�mDӍ��B]e�3�oj�t�:�p�{����!|>���Z}IfF [C��=��8P��5ԧ)����*�^�hKU�<�� �2+���PT�S�h�ۘ�g���c���zN6��J����ah�P�@(0�B����g�d{�HJ:����d���#HX��H�T�cL�r[���`'`���Դ�*~MWs�mu4�m����3@�O��CZ
��^4��q��[�#Mj�֗�RM�z1rt}���C�����y@�TP^�����;O��a]<��Ry7 ���Fi���ާ��	v�FW4m7�m�$��zg��.ȍ��S�E\�D:�}�pV_�,2R��L�t%eB�!�~��$*���FW��!@���^j o�a���q�w=Q+�����N}�at�q�� �SH�g1&�M�r�w
oq�����V*bD�%�Em�R�km�Ѡ6Jj�RJ�v��_m,ղ�E�`���6�^�H���V�s��ңr; ��GU� E��0- Z+#hky�}�|L&��/�pP�����Ai�)�T%�2���i�)ґ��B+�O-���|]L$ζ��e0cw��F����_�RlK��2^��6MeI��q�8h߅��b0a;������7��m�Su����Aw�7�'��B��.Ixk`W9�"7.P]���F�H���ze�v�(��]Koq��@�P6Oz�j�Kk/MX �ۊ��
�O~Y_{fs"�����H��m%��\	k�L��d^h��s���PG��Z�v	�H*�����_�Օm����y�[��k�v�����泥/i0�(���p���,">�z��7��ɖ�;�ƊD=0K�:.����a_z����V77����sUm<#u�Ƽ��,]�/��UT��C��4=��V)��F�ٜ�F��*Lנ�d|� e���#&����`��?L�	��`�"���H�U�}��{Uzt��zz�`�:+&d"�W��]{bFF_�4ず�T|��9�hp�t�a]���$�xgSp�9(�TMqɦ�[�s�J,�	�=��#�MI�؝�s����/*g>��{fҼ34%s*��2���~[�]\�I���"����^��O�X��q��e��7���LBie��8`T���Jt(�?�{!��?�V��������j� S"� ��~>�lq>�)f�=�����"ꏦ�V�8��UJa���6YOy��{�]��ճ��Jo�'�S��E��HX�Y���$+���8%]���p0��X"כ�-e���1Q�T��(Ѷ?�y�$�군1%�z�`��p�����:��H\g� ���8�X���Tڟ�@y2�@�U��?�,��-)�����l��8��h�%� x���m��u4Y[zu4.���� ���be +,4��/��YZq��џ�=���8����v}8�[ի1�Y���6:�v���e��ع�pLZ�I��/6y��qٕ�=���+�%!��cL-&�E�|M�F-K��CN
����	���c=@'���dWN�VTaH�9%t�_S�����S0�^I���U7{+le⫻?5#^�Z���[M�$èl����oI�UR����-V�[Mf`ῴ\m	�Tbf4��o���`�0�����6�NJd9]/*+p�*䎙/���%��@_�mEz^��V���R�u���1v�tP�U�6g+ǋ;z�?�MD��Y�J��d��hbxd�K y�ȣ�#��5�7��V��U�PV��/9�}5?��p���(c�ė��ɐ�p��1NG�n����(P�kB��:�]DХ����n��f%AgB)8+I�z�%gh�a��\���abn=n��dv���[�.v���hWp.�j[��$�C����׆��Y;"�~��揩,l��i����=lY�׵{5��;�saTl�CQ�Pi���[�������B���~І|61%�^k3]�RhY�h�縀v�/Rh����Uv�;z;'��s�ur��!
Ѵ�NH��SoE�Q���Ed�)k*�b�B��7�_����wG�R�|G��8ˢ.�H��FS�
�@�.,�j��,¡o���e
�9W���D��f2Z��������}ί �O�'<0�}��y���Q;�)?�!�$7F�g��Px�7Ձ��j���@]��`�%I�
>$k�L3R���'x�'��������SY�o���[�01-�~+K���y�:{$T��-����'䜓���\��DU���ү�1L����7�����z�r��~N�SQ �7�s2_���cV��B��&����;#�0�e���~�O�Йќ�c��"�֜��j%���B�����vs(���KE{���2�s����$/��EZ��ɡ�B���V�ev�����7�=�YÛF��rf�CE ԀgG�UN����2�ί9<
G�u�%qՀ�E5��^d�f�M�RK����x$�;��u���<z�$g�vb�׺G�7;aB[���%�J�q�l�w�1U�;�Uψg^eu(Ch��*}�i�;1��c�t�;�TEiq0Z(T���yʁ��sƹd|3N6@ֆ
p"�s�HُY�M�a�䇻�#q�0[��(ْ�M��+��c7��/>40��Ҥ�b��AzW_��I.�*�÷�
cb�@��O��#�M�
�wH��N֞7Q�_ӷ�d�٪ϕ�X� �1[����s�����3�DL�j�F0ƒg) ��@˂�\���Z�3s�?� ��ʂ�q]���f;@R���*&t�d@��$濹�F. u�A����g�O��w�vow�"�i��5��!�#S5���IQ�ʹ;or�bc/�ٞ�jV��z� ���;_�����xyt+��Q��sVE����t����@���=g\p���E��\ ���n�2�3�$�6�g���7/���B��j�t��Q�-�:IbѤ����J���([��<S���)�p�r��*R�E��"n�� u(�T 3���RC�§�#���|��5(')��)�+�&ܺ�'���R��Ny�ѓZ߼��Z�b|���:è��癠�ʷ�r��f� ������\{
�7�1���y=x���ػdl��B6S�VP���"F2�H%c��%Řf���Y6��{S)����[CUi%T���:��þ��"2s���1	s��G�	y���ƍgP/��� �OYyUh�K�da��U(��[�˼��{�O�Ӂ��p�o����%\;z���c<�%a^�s7w� G� ��e����b$�!c<��5��x�S��=�c-h��6�XM9&t�"]�^(�]�PPܥ���%�8�3�"x ��l����6!��t�4�d�aK�K"/^��Ť�T�_�=م=�IF�iԒ����+����G�hI��s�[5���}�����GǦ����W%'l�@���9_^���x�SUld��k�L4����{^��/�S(Cey����W�T�D�\Sa����K�t��)��<uHn� ��R�h��p~����G����Mj�
ht��)b3�[m/V�zF�U������׻>C�֍�h�Y�8�%YsU(1�=�'����TRWX(4'�Tȹ����i(��c���N�ƴ	��g��=Ec���ID����O���KN�J�r<:�ڟy�}1��`�x������kV<]	fw�An��@S�Q���Fq�IdYľ���.|���j�˸Ə;���W������dm�����5^��~�+fѳ&'5O��e]x�6k��W7`�I��$U�a;4���;�=w��~��n�}!��O�yx�
3a!�P���p��޹�lL��*h��;W?�����nR)2h�/c��&̰}�?S�+���B�{���ɣM�n��雔��y�1��׊r^�7�]�e�]ЯJ�M��O���|����˳A�7��4|��y�8�
oˇ�z����bIl��y26�g����K���m��l��aYH����,��I���$7��N��cxC"br���>ߣ��Z���Sd"[�@D�a��u���g�ӄ���Ѯ�'�a�v����Zi�&��s����j�z���!͈�Z��}�/������*�cw�M������*�l�g����h�C����v��|�/�c��Z(���;	�����ʲ�2QMϣ�s<�[��{.@�@�?�� �J�����"q�]�v���|()�w�+#t	��d:�:Vf5��6����<@P��n�n��
�1���Q��VU/�������]1��GPq��j��Zv�˼�p)�>���.��ZC�_�ը�&�'�T���f-.E�Ԡ
�l$Z�CB�~2Z����(~��k��5~s��݄��q�#��fʷ�@MS��Ղ���4nLSM_����n�w���	�&DP����g�m(�]�@�:݋CT-�2�U��ɛ�(����"z[����i��u:-�O��������Km��Z�[X~�0qkoa��ه2�>�{��i�O4�۽Jܳ��װ��l�,���־���Xp=
�[ �}��yŞ��Tch���mh�Uz�Y�`M?�O�k5O��㩦p��y�?�H��Yo$�F�>2b��DG+���,�L���Vz7N���	�g����׸��&:�
�Y���^��E$�)z��y�y�Z��td�x8L'�j��~�(V6�K�GU�h�~X���#��$\uƜ���$ݤ�3�l-�
�
��kHĔ,F~=��*�fV��3�ӛ�V�/�J1|^� rVX��s'��%v��d�#�,M���_
I�a�7����Z�8-	�@3\F��YuVCN�]��XK!�*յ���^��� :Z�a�m��Tt�5Zɴ�����#2a�[?V��W�zDs<=����ׁ���D�`/�v�$/׳���e)���b�M���t�JDZ��[N۫�:6���������^���2עs�	"|h�e y�&"��j�6S��/�L}�	�Kr�񞼯�V�ř����Қ�7I˔/�-3�K�dU�Ԯ�3�����
>��C�۩%ZvU��\�"��d��5����Oi���j1;_���Lg�
gW[�p`-i+i�v����#S"n�{�G+*�p���c�!jJ�3뺋�G���=z	Ә��,ͯP#}�oK!��Q9�-)�=Qlk׹
E�!���`������a������D-�D�MT%��'�=�+��}�F=�٧����'��RI�	s��>�<�����Lc���`թu�D[�k���J,��Bj��&ͮ�\�>�a�:���=���Po��s��wJ'����B�'6�z\XUC|�oo��)��"�T�Vc^�7c]���.�}D�m��i'�2(?]��b``����h��Q �mwr%yoU��w���,Т!l9��7{�ݐ��:��lF�9��|�,�Y��A��H9į��lYy��ݲ���hO�
.lI��@�R��ȼ��p`�Gɿ]!±;����oyV��߽#;�>�C��V����I��/���)JM�B$%MMfmV<���p2eo ��)�f�S��^Х줳����#/	�'
��d{[��ץ�ځ-�o�׍I��C�l�Hb^lBӷ�7yM�qY�������r"���c���[c����5Ⓢ��|�0am��5��8��%+O.���_��Wf#�Ư|db�[v�&
*�����"Q�:�8*n)���qj����Llx���h��|�B��%.��P9 u1�����|/`]]'{��8 ������([�#���O������(�Uܤ��v����$��5��뉮8�AJ���WZxPk�q��j��!�E�\Fɍ��Κ���P��\QBFH��>�X�-|R~�/���ч`�ͥ5E�����7J�i4P�qJ�@���e�d�'��T�oͱ�^<����| �L뉏 Z"�R=�{;s�$��
��%��P.#~"E�b���!L�I��¿��dKڤ�F@�+£��2^�P_��� G����×�/Y��#?�ݪ4h���4�0�o�KC�4�
q~�[��-����I�����*���<k��^�' ��uB�g?���f�w1�����n6���,�6_���D}��lCA�²�^�GnP[%E� ���LP������;�����kz�"l^��^��e;�����D�#'_�A����of������� �<e[%f�>>�4~Bo�"�2��,rB8��9�.u�N���JLaw�6꿐�%�`ɩ�QI��	
2B���ӓ!@@LJ���Ɗ�2	ac���|X0 O*|�W��O&�x�#��6vg���=��9�b��@'���P���c9L���|��*���������y��	�+� �22���� ޢX��F}X�U[e*_6�ԕk'FFl��bG.�gt���ڏQ��w�%������+}A�����7���P׋����̛=�Yf\7R� V�v�A��S��f,Ѥ;֎�j-P�C�c���tS�w�d�y�W*��ϑ��$��m��Gz�3����miF��3AJ�í��q`�0a��JA���:�'`~;�P=�}�����γ *9��pn��q�W63�1;|���#/l�i��J�J��酶��c��Bxnn���Jm(|�=@�0,g|Hq<LV��Nj���Ns�e]�u�	Fp���a��I�J��zPm������k��КE������I>l}���G�4�_=�"3�X�b�	S��g��pq�����&u����f�ʽ�I��*W�(��G�]aϴ���Ɲ��U#섁���׹l(�v��~*3*��V#o\�_Ŷ���G�렙#~���$���&�������>��3�]�#R�o�x���쐷�ǲ�M���B2���۔��"�/KfM�,2��dv|��E���K	�{YpM�KJ6D~[��C�������m~s��I�)��X��7�����]�3p"�4����0lUuU�F�v�,XϨ���m{dmtP˛����u���h���T�X�N�r�1������1��,"KD�DgL�Ï��H�\8gP�OT�:��Y��k�40��ʘLR��ņ�	�ji'��.d�d�E��Ti�Km��gUs[���/�WR�*�a��װFQ})�c��g~�z ��{�wb���Z.|�<������Z��D)n$<$�żaE1-��矺T3G�a�jQ�{��]�G*$A9`&~Z�K�}�]x��+0�U
���3A~8j��6��}�O�ܑm�"�D'�{K�;�d�(���.������m�zClt�]���X�@�j�!�'���K�{�w�f�`���?Vmůg!����(��	�I���PKA n�!xa��|�F&�$K�$֗�jY�⼝��A��ϯ"6e�;�f�-n��w�_�Ѵ�G�0*v���K:�,R��E�Fz�D��=l�zI6�;�/=��%|}�[�K�[�MK���cK�;qn��^��ď+�*�vqB���3���{"����#�&�x8��3�14� �>x!�6D���e$���zu����D��I�K��Mj.�`U�J=�L{a3˶��NS�����n�������т��,]W7����\'���c��ZP�\Mޓ���Xt�X	�w�_�/�SOPR����^����D�s�Ŗ�����u��I6�`R^d�������a�m�����Q��qci@3�_ˡ��r�yx2�R��f��jv1�K�4�5₣�(�"xR�<�D�Vk����p�����ᨾ�8����nk�,j�^&˻
��[����uK�.?�?�/�U�I�L�Tĭ��d�U~_S��&�+ݚ2�62;�ْ:�A����4�#l����o�<G�o���g�#)+���iZ��eZ|��c"�G�����quv�[�`F�%������ܱ)3y]��H�V�ٙh#.�F��Ȫ��^iu����ЄtK��B���"_N�ꭓ�VP�XvF���e����Y܊$a_F+Y���]��ĸ=��q�J�3�c��gJtr���o%�^T��~Y��GQwv����K���Cц�X&�@Ѭ�سr�	���g���j�B1��^:t5�>r7g�<�X���tήܗ�Su���B���c=W
>��)���8	 ����^�D����4u"��b��s��9�jJ��9e�A����cV�P���TUz�R����_~M��_KÜ�_p��XL�W�������]��ة�aTz�CP�
�_��[��F�M�b�ݖ{��y��[.�k
�����󺶖;B�YO��*T�Y���4���)V��_��lޔ",z��)t��Cn��c�����Ml�S�E�=ќӒO�xU��M��b"4��e�`�zo�\Xck�	���
���4[;۾},`/���z�H�h�6�/��$���W���u�T{��j��<xD�O�4"���u�/��x�Hu��m��W�*zF���tp�|l>���j_��i�^�&�i򧺝����_I�B�<ĵzL�~�f�< �/���Pf8yKi�8����qg�DP�.�/�1t�e��J�O2鲏���&��ra��S&4�M�I~nF���t�܏� �Y1���e$"�����k�����ZoHo��6�!�Qe��G�w*YܴV��x��wn�T+��i!��Gl�������T���櫵;�^�&��QW%Ҋ(����2���Y�$B�������O5�O���6���gJ���WXr2;c:�"�Q�h���9��r��a������j���T���}}�֨�QR�d�27*�'K���_p)����~�/ :V�:9���Î��X��3�ꛬ�I<��?�rе��Z�����/"F)����6b�T��  ���>ϰ, A��!O6��׆�U*�1^mBH}�qZl>*�1��X��~�k=�������b_�d&�����Z{���ڔb��c<�}1ي+��S�y��j�[L�O�6���~&�W��	�� ��G�ǁ- �X��1YCbN��e�~C��?"T�'�.,�3<tf�14×>�l)��g^&�l��J�ޘwe?����y��V��NN�h����%#��������
�ўq��v.0�%�c������M�Q�O��S1���L�Tۓ��Y>����Hg��h�n�@�w�,��94>a���8ڥF@��jVأ��G9<oJK/u��s��,2�ٌ�K�%)ſ�%T���1��I{;{R�@�-jE��O��+�r?�,ک5�n.x�9��g*��px�y���ڨN=��e}�)���좈)�~�]��T�7-W�����*JP��}��r�,��{c����_�����#{��x)�=��]5�_;Pg�-���~r��ǟ�HޘM�] $����ob�ucI9[�Bf��MH<.8 -X�Ψu�/7@p+�<!GĔ�� ��u�/���* *O]�6�Sh0�w�7��]EM�7Uu��|���2�Y"�DeJ�F)��v�Uw.-�ؽW8�0���� OLNp�ٛ�jt��T[��j��+�M���.��$��Te��t#&���ֳ6��� �� �&������������>dB�@�L�C�w_z႗����p��|�B���<�=�=R#��(v-����o����4"|�:�pv�ζ�aH�6 �װ��Z���M3�V��j�1�D�k�F	�Il2	VD��<�!,  ��=�C��Oh��~D���o�ëE{�m�T�@:�t�Ԉ��].�MiC
�m���g�/w�LɾF�A� �	��z���J� �����{��P�`��x�ը�U
��Wg[b���ډj-LM*��a\��Q0�SQA���������L?��{\#F- mCd9� #v$���4[i1�V���n��R�A�q�ź /��j�đ'�o܏���2�ڽ���9�a�nƆ��;��6L9��X��׬5�	vv���L�X��~fh1���6�o[����4�L����p@{����WR<��������4�V����\����L����m�{����z��վ��8c`䍯e,.t�1��$
j��(w���*��Z�3} 'T�8�5(���Q�>N�)F�~���,�oI��v�ש ��P�3��6:57=SH��~xw�O�w�2_@_ e�
Œ������{��S�.�7%$�A��˝����@נ���,����P[�%JA���%�H��K9��?0�[DO�E>��q� �e��2�^�y|�B"�	Q=�H��Fr�V`z����������c�V�%��A�4xxjXEE�&��}�n�uO[pX�ѥٗY�FE�
�aSnOG#��hS'98_V�N:��r��FT�@�s�R�cF A���t����7��=C Ϳ�%��W�"Pm[l�J�2���;ʨ�Dw�!��w�,-�o�P�KYf	���OY���6{�^��7�D��u�"W����@=��@�C�bT��g1�B����*��|�tt��s�j�|��F�>*d���z�� Eǯ��}M .^Q`q�`lf�������e�UVps��Do�{w�6NF�&���2��m+s�j#��X>�'�YQ������r�ѣ ���j��KR�m�g�:�~�ٔ�.����@��s1��6�RI�{��?&�k^{�$�����>>ĝN� �*���u��%4ջ��Y	��8�bP����hԋZ�W�_�G�O�9�E��"�o=��4=��^.D�Ê_BEGN�$ټ�꽪S���8�2���ک�$)Yȥ�b��b�_��,�&�	Jk�{½�Rq�S:���I<	fV�Zp�*�<��('�0��T$������I4Uf�>ĺ�1*=���b��+��t�B0�'6�tX��'�2��?�H��=�n^Y2�/&�<��)�9���n)����TK�e	�p�g{;�P�G7�̫Pbē>\�M��������A��|�,䰍�Ĉ��89
y�:��o\�,�B��h��(�
�&�w:��3����TNT�C9������Alŀ7�S`=P��"*ȒD�X��p�r�c-�I��W���N��j^8S�A5�I��*NyJ�����-�S୚!��v�Al,S��Ӕ�� �����P��+�e�!t�d��@���U����io�l;|#Z�P�x��P1��7 �'dc\S[�\�ը�ڹ���� ���?�M^�v���r�'�|m�ԓ�����:\�ʟ!S{n���B,��Xy[���o��d�Y��5����y����o�%�R?08�n�*NƈY�@3DR�����0��m���e5@��ɤB��<،��Q�����!�̝������Y�}c�#]��2F)#��q��r]-����(���?�#�?���C
lqáGz���ڙ�B���Qh&�^l-i�_�)�B+�����~�=r����@���W�B��V��{�:$5Vh�JN]��݃R9�;�A�'*�clC]�z���� �����oE�[��µV�`�&�BVT#a���I���O��qH*H�YwA���ͰE��N��_�X�f{e��B�����8[�9	ф�}���	�Mp�ԏJ�z�h`3���ap��|4