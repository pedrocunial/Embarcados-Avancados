��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c���ѢǓ2�Su���;���L�X��2{�ԑ�(I�lR����+;,��ؘ�~giאP�Iq+�	�!��s[k��h������HC��#���W.��VH��m]�Є 0j�]&���E=*�A�?�My������NC>MKw�2�5�p�M�P'�|+w��F��i�� �����_���rz����V�����"fR�֋ԟI �h�����5��(��๣����yl��8�1	�&c��$*���>6�x�!���,��9 <��ފ��Y����J�|@�钡#|���x����o������� ��N[�T��ԝV�sll���>���B�h�����aλ*�D9��Nt�M�=bz��i�@���Y�֜��RQ�6�����,,x�0Fo��o#9������0x�ʁ��IFF3��">�� u���ԇ�ә��I�Glp����,�?�ך�_�15٫�gED:,���,�q@m�<j��w�S͵(�v�e~���S�+�{�E�g]�¨��ӷg��t|��ԃr�9ys�H�NV�v},�(g���Y/ ������6��É�]�4�+ �tU،�A���Hz�$eq%��c��a� 'f -� ��F��L�\�'Q�f�Y�r$�i>�H�V��؞��у'�@��6{�)`{���\5X
Cr�a��
���O��0��ϏH�{�j40��A��k�YW(ƣ��D��yC���u���z@[#�����/;z���KJ����NF
R��p?�����&`�ACP�5�3HLv��RW9�hA:��H�ސ��yK	0�E�kx7��Y���<�Hp)�囒_В��(�~�����JK~xUS��;�4T�J�279��{��SjH�սal�:�f����h�W��rМ�[8@�g�=�)Y�L�`��u�1>����CN�TRi�ċ)&.iwM]sR�a�9���o%efy.�����mc�h����7�Dq�,2�S�<�u :ҩ���D�
KCV����{	U�*��VQK�q��)`Tv�p
�����QsX�/��j��l�ʝR<���bJ�dkd='�5��8��Z%�fFR�#�4�΅3�����I�k
�l�M���N���h����ؖX����LȀ�i_5�N� �uB�������(E�(x���h!���Ş�EB�� s�B%�a��L~Q���][�+%F��6�omV�D�֞脦�T6;t1��a,��@%KX���KU�zPl��Ɨ��>���$:
ޖ���.�<V2�R�(q��E&c F��X��	<�9����@�1�����A�1��@�v]���	s%0��׌�3a��c�Ƽ��Nn2��y�p9���
�E"���E s��i��P��)0��uW��+���C�İ"�;
T�aQ�*b���3=�eyW\B����
GSGş��>0��?:9���f�E!ȏ�����_��с55�Ʒ2�UCU�G����%�����(���0OP�!��h>҆��`��{�KJ$B���&�D�M��w��z���Yby^[���i�}1�{T�Elr&�;�Q��_�^G�x�I�oǫY�~����7��U�r���zW�+�Z�\7��U�<�.b�8���`X�:\��Cr�绔�TK�t��ٺl��n�����,qj6�IWQ�j���7�˲�?��&�N��}"kK�8�.�
vZ_Hc�r��K;����U�*f�6�
�%�����
�����êv�`���_!�V�M�LI�6��6���C����!P�R+�w��{����|3��o{��1�\͑��E_���5eS�������I���R	��G�m���� ������ݞJ���M��;Q5�up.�oW���۬�r�RתE�EJ�7���ɠ���W
n��n0��=&��#��(���W��`T�4Ч���i=�����&��x��2�����9_�X��*���|;�2�x��i��R/�M#��d�Y���B,���td���Ol�+Ga:{���9]�S��C��jL��6�;>��4�Ǐ�T��.@���
o.E'���8�p ��Xt֤#��B�\�;v}84����k��7f��)���=N��(܈�r� �����Q'�3GҜ�-?Y���_�:Y����q�:ر�R�����Q�����uwK�2*�����eI��.c�����UC|'^�u�%�$�+����Fv����o�ϒG{�W�j�у�o���V�":]k���F��!�v��9Nr�������EJ�цe�Cܭ��U��	�X���<�X���l�>�����mf'����n���厤>������S$A���k�:�P16��,{	'y,�YO��)���m�O�u�[�4���O�Qf_�Mm��z�J�����=s'���V��럘���\�w�&[���/52��	��rJ���K�1����j�����4wa��Y�ٳ_��]�k�\zh�1�*r���'�R�x�#ma���<� Б��a\t�̝ΐ�玷�`��5�mԖo��ө��߆�d<��+Z�pԺ*�)�c7�Dl����r�!��ڢ���w3�iͯ�j�K ���ێ� X{p���uyD<��9v�担`�+��@໌��Ȫ9tݎ�Q�;���i��G'N�c�;��-�:�T��RB=��P�e>��1H�e�Τ�<��wQd��Z]{��.���[T�4ժ4鿷ѩdc���"D6ly��?��4"��e��M�yt7��s�ؙ���wK�~<ų��7��o�����j���Q'���eҢaB�n�8���F�� ����Q+�\��?�2b�#���r��y�V!�酨�ͪid��([Z���t��{�$�"`�������TF�Ez���O�������"�yG�l(X4���(�����sƖ�q}H�O�J AWԻ�͌'�K��J���
�����l}h�������%�N�hS������ #��t���i�Kתփ���X��pX(�%�F�::��;|{��e?�!A��L���Γh�l�!T�aruF��1[y��.���$H�Uvs���MW�-ի[fN�W��H'��V���9��u_�2R�t)@i�;�ג��o!��ڊGy�ӟ�{���[^�뺢���8�h�a��'I�K�]7��]�_�H�"EH�b+�0���f^<�ˁ�T�0Fm�z��.�����Ok{���i��	1Ո�V���q���G���w��O;�HD�x%r%B��XrKv��8[-�љu�a]Ü� ��Շ�iV�f����~�NJ�k]e&0�[΂�z4U9ܜc�I9ۘ�@$����(EfQ_��Y����	��E��ڍ�1Q2Q9��'�%v�w}�Y���}�'��1GL���-��P��� ��4 �D{~0J�Ea�r+5��-������$�y���^M�;�w��Ϫu�",Mǩ���h����h�TXѾ�Ѭ��>��?c2j=����?��\bw�g��bP=E�j-yM��������;+��w���	�M�Z�Yq&k���g����otY��۾��".�zH{���^�Ա��E�.l_���#� #^��ۡ��;"4�ȅ��C��5�HMX�Mʡ���E���A��l��o㚇�_�V�N����HƂ �<5R�c���#j��R3����a�q)P��M
T���B�}�F�(d5��� �0x{���̮�9����I�ɽ�mè��fZ�}��6��LnJ��[غ�N����� �cC������L��8� xwb:��-P�V��cz���h�ͪ����C�j@�2L�wY�8�peTG{�=��h0ɉ�K�� c�)�`���P�J��
Mݽ�6�0;(ZD���J�Rl݌*iQ]]W-u�Vcv�Mf�0HQ�3I꠬����]��vjU)�d<r+R؋_&��`Ƨ�OjqT�}���"�j1�1ZFK��{"$Q�ʚ=�}D�+��Z`�Ч�&莳@�z֫l�d�35.-�r5��7�]���Ah�E�Vu�ׁ=�ܰ�^��츝нp���Ğ���d��rI��P�Q���
��sN5	��?5��B3��l%YHҳ�"r=!�# �h�ur&y*�������\�2����?��w���b�!�橠�q��ٌ3\F Ω��R�Sp�ϼÇ��$kdkA2s�j͏-�bL�^�}�P����}hL�� ��B���J5��$��ť��U��~�?�|�2Y�1Ғ����W�9-F�m�z�B�l2�>/��"� �4�r14���4�R�[����T֦f
��vx�'�c��	�E��Ql�Y�G$j�|¼:��X�ڢUߟ�i%dz�-^%;�k\d�3�F�;	j���u^{�ı+Fx������ �?��h��{MS1�����(Q��C���dRU����@{2���a�d�ph��_��`���c?���l���.4N����1�qT�tp�Zr(p�Ff��ef-��d6V1����k����h�{����o���<�Ήd��U���6[w%��k!��8MQ�9' �*��oe&1l�N}� ~� ��o����T���8BBȉt	,^��Wn@�.�i�P�XO����kl�{?"��������*�,���Jf���������/�/V�����wW��i�@����o5&t#:�n�
��fGT#�����ȶ����v�� 	�r`�P��e�����4̹�a��d^�����I�"��B#^�+������
KJ)����6�Tg_PM�R]�|�<+F��%��%P@�1�l�';���@CL��o�)Ԧ]�����wѮ��-�����Y|�^/2��dΓꥂk�-%�yp�:�b!X�I�b�h�W�3�ՙ�~���S+$�FXV�ckĒs����0-�{�:�������U�29�C��=w��6��]�-��C>a�G٣�͸�{�gvf=;@��td��u@��^��?ҿ��!k����W�ɮ����3��B6��y��y�w��ia�r�+UxԐ�<z����,W���M�Ξ�
��b&�|�?R
QwCm�좛E�~D�TM`�(	�13�_���`l=�������ʍ��s̑{l�a���V�d�ת\�<�����n^� �̯��͛�.����b�$����W��қޠ+�=�H�.m+)��I�@!�t���r����i�iz���2B���.p�@�_�[�MC�n��Cs��fz��H��T^���C;�D#��J� �JH��lf��пLG����m
_��v��sm�����S�v(H�LCc�@��M�d��{�V�"�^��l�3wXkSH$M<v��n�:Dv�6N�*`����I�=ɒ��;��|!��Y��,T�eV*A-�X $P�6�^�X�ш�50\������)�^v|�⨻X��i@��bD-J�<�!f���:#l{�gl�H�i�ǟ��W>�rhR`�$�*�������*hS&\!D=N3��2��֬�P��Jq�y���B�5[U����Is�Kmc�-%?�����SUm�� 2�\D�PJ��܍��}]`X\Nz�b,��2�r4<�蝾+�;x�\�5�Z�6b�MZ-��l�^9�Zk!����#/�
��>��+$��1��!����u$ ���ѿ	�(��.핸<<L^X���[v�������������Dߜ\M�g�'��?��C����6�u4r^Yv����豝^��;���B~��I�|L�{�j�F�ב�F? �f�n+���L���(�M譛Ơ�,=�u3Dz�z!D�F��Ei�NT���t��N�J>��o?�ְO&n�,����\��r�w1��Ԟ��,����C���O��x=mT���� ��\R)*�Oꬖ� WXB����j�;�'��z�t�͇w� Yy�,��Mt�iܿL��y��,���}UQ7���Du�)_8���!�=�6iԉaxh=�"|U�w@�J^�H�������۽��S�ƛF(����<]C#�N��z����De��ܢ��&t%���ȯ*-���! �5��*��l���8�L�[���/L%T����X��.aL��a�BI))fbS�e�F�+5JOq��ڜ� ?�%`�(�������o��u�ަ���X�yI��9�HC@O�G�i�4@�uH40%I��
�ι�3�f�@�Ѯ*W�kk4�(���/����M	k9+L�ƍL����/O��[e����M���t{zQ��_P��B��~�_ܔԾp��)��������%`�_�����#�~��@1����ph�!�u�=%��O��ܴu��&'`s+��|5������Q�R��"�z�-�讶����[�?*��Q-�;l�槌��ƼN�cu����/8EH~pG4)��rD��K�9hX�xF�����M��fUaի�곺�9V�5Ɍa������B<���e�["�L҈J��"#�����Q`��F0�k�A��4L��!:���v߶v���0na"��<w-��f�����АL�C����D���X�ZFɲ5���?5��4)���x�D����ٮ�0.SO�r:�u��`J�=���F���943�{v?�sk�p=0)��U#��R$)�< �&i�<	|v�1ɝ���o�j]'1�$�;ٚ�<���Z�0C7����$�8�`��ǻ��K�i�y��5M	�dى�cS�J��uzX��G~�ﱫ�-U�$���������ȁ��z��l�����t��A�Y��3���z�j]+&���j�f�-�fw�)���͓&ݜ�ץ�{>M[v�jY�;GQ���G�W�˹���o���cM�����F�ދ�PH���~�?'�¶7�B�y��,��о�D*�����vk�@�oL���?-�і�� �$����*�|��T�cn���D�	a*�5�B���[^{�c:���+�ԦZ�Z�Ԑ���s��Nu}WJnNB��!OG2}���r{0��s�\e�`�Nl]��);&�5y��;��m�i�{�����P18�O�.w\ܩ������ lXl��ω���3�����m��|��~�]ճϫq�b�]q�-�+}�3A)n˃0Wl�(N'As�e���Df�\��v<"����X�DT1�i��	h��ք�V6(O����|I���o_�]��+2���7�����9��'�>y�[�VY�g5R\XFq�@�e���;ͽ��~��_M6ŧ$G�pN=A7��;#�r��Ҟ���>#�7�蛲��X�v{��Q�2��Nu�żם�jX�rU��YݍW֔���FCz�gsL�e��G*2��{]�5���E�^�,*́z���-fBb3j�H���;y�2��N�4{߆TʏC��s~�s��~º���Z���\E|ȕ`
�9�;����ԉrc/���C1���F��ֿ���8��6?&U�C�}���!J��v 6!53��f�e���o��W<d[WZ�'�t��t�p[fO��`R�1�\��9�!k�eߨ)�1�G��(8��g�ގ�$Zx7��,_7{UK*W{X`�H\V$�Z�l ��0����.��f��!N��ѝ0i&��,�K�f��fe�z��?�{��\��lL��D�R��q?b�)�Jҳ���&i�sƷ�?�Z����Ǟ+ݹ�7KϻR��Ӎ�i�.-pp�z@�N���S�U�MPs�j���AGB�<d��:��I8��4V9cWd�?HP�g�L��.��\��I���6�J
*�?�n�	���12��=�E~���4���ܕ�.u�����e��1�o�����M��+6�9���+"���{�����/��R�rȤ�h��_1�wfU�4N��1�R��%��q��4}"e�}cQYW��&�a�E^���S,�g"��#�C��z�Q�ݯ"���{���8�K�a��0vRt��$d��qذ8�aOh9�j��F�j)v������qƻc4B-���:/#/Pǻ���~l�f��r����#��E����a-�
��7�7'�{�&�B�
VS��E%B�*�J��-
�n5i�j%S�����`�p�F���g�sT��)Ӫ�7Ю���(&�G%�}�>��8MC�H�q~�`g.3�*������?�l`.�F��(Te��&o[+��ԌpV5�Tfc�3� a� �1��Q�Dg*5����v��Ә"P� �{_Bc2��E~[��.���<����� �O��
����<��X����0k{��H�Q�v�M�e�fBE-'�)��f�KF���J���w����#:sl�-@+=�RZp8׌^���y�
�fN*b{2IJV��t313��� @�XT��zC��kiDa�>�9��d��?q�/�\�%�?��p-yI2�����0-��5rÿ~m"g�HD#�4���+�/eg%����S��������-qv���)���֍�����	j�j�;��)n�N�Ba݄��c�q������Y���l����6�,	�Ȳmƃ���C~g|/^l�p�� �Ⱦ��-�7'��,�Ř���7צsԭǴ����]7���Gc�@e���@�g���fU@6�.	��]�_�L
�ߵ��}�>z�R�Hڞ�g���� �2�!?#��ާH(��X�J�)�15��j��'/�s���p8�ɋ��%�U
�U�a����J��ն<�?�وg�=t!������X6֌0������7�ic4֡�4��ATO��DO�r��_!/6�����?s��&����Rd����>T�僅�u�H8�b/PI��t��T�ԵѴ���YF�������Ϟ����)8G�4[��J������8�n^�6w�+�[���p��?�һx�	;BQ0�=<>�k�|��^�O�zg�F��~���0�Zi�Ń�6ěib:���݉��OAY���%}z���[6xQ�x˜YK��p�`(�3`���������N���=�"+��P|߂�;��Mċv"�x`?�jK���֔���x�n��WIɕ����!7n�G/p$҈z&�N{:|G�⦘/��ӹ���QS'"����x���Ӕ�w�Y0�_zE_��<?�7���5�rg�VA?4���x��;W����ɕ�H{�"޸H4��Jy���hIB��)H����m9e��D}��d�yM�ņ��h�6:[ڭ���d���7]����穞�h��U��WR��R(��+�0;	n� n��Փ�va�a�r>;�n�erӝYq1�l��Oa2�"q�4l>��D���1�hU_���I���<|ZU�?���+D�Dw�W��*���L[�&0��lN���S���GK��=J�B6�49�ɸ���R��-]��KJ���1$:�,�,o��0b�{:I�v5݉*�-�����p�~�R*d�GEg\�x��H�4E���327�ٶp���#<�||�bI�%�R2f��l�5ۥb��^�uȒ�Q��b�E��3��O+G�/X �h��л�6lC/r����@�V�Ӌ�˜�
���{eN��։����щN|C'3N���âW�o��J������O2�t �Ŀ�����h��M𱇋��}U|�?��Jt��w�:\MyM�-ͤm���pTL6l+:�@P�]�=��	��3dn_�x�v�|���Ro���~U��!�;�]��Ϯ���GnS����X��U�W�x1���h�]y9Sp3�߿��`,H�|����Rv��	�I��<�= �7Wg4�����G�:��Gن �髨_կ�@gfd�חX���]R��I�J���^���G7�r�	c���H$P�Gz�h}�#.�K����3 ˽�9<X ajso"JR=�[��e�B��� Tg��:ׇ'e���Wɗ%�m<�P��h�iv.ERqg_��ɃҤ��oYa*[������}�7�G�c�}��I�f�Ê���#�����D�m�N]��B�� �:H��yn��/���n�c�{�u��ڟo?�ϊ���㚠���	�yK��#�&�`�$'LbMEQ-Г�;**�ε�����=���-�7�_'f���~�¤��5i���{����2J�+���Yȏ)�Xsk~'���G��li➦�k���(�`�/#���e�E45#f�@e;:�%}r�����xs���G3��o���䒗Q�
�����*H��?��C$��Zo��u��� >^�-�H�;:.x�W`��t5���j6�К��K�z�	lD�z����Hy|�!��&��ΐ1�r�8�t��2�6TRM��ߒ9ZN�X�ƺI����p��ˀb_!`X�ȃ�})�	A�d:��7�M
�U�^بN�+u��a�KS]�Oq�� 6�`�N���1����VxAڌ��3!D�)[��ք�~�^H�i7����ε�~�c!5���j0Xb?S�?��@MF���>��������z���B�w����P����?�A
�70Z�5u�<Y��b�l7}��~��]Pt�UO�"�R�v��@4�r��L& _�Y�V��܈ۆ"� ���kjy���C�N�L���K�=����ۆW���o<ր�����ɍ�e���Ӳ�F..���~e�k�F�rv�#�^�&����װ�OժLOuHvW.8��݄�7�17�$.�N���O�q��4�*g��꾓f�(�f.�Z|��@B�Tә��>��K\Dg����� nv���, M��t c@0�B���a��ϒ��Q[$b�0la�Mt3L$�怰��S�{s9�=I/�߃��>��D��8��we���P'o���}����Y���	�SE6r.����G�Z�8����4�Q-s�C�K�o��mی\����ح�� ��N������tI�u:�GT��~�|7d�C9�1��8���lx�(�d�НQ��K�vH�"DPu����/��捝�,��e Z��������{����V�I�-0�KVպ�2���h�Q��M��oh����Τ�q�j���v�`"�Z������K�i$�d���A����IMQɉ����}(׉��<�������o���h�K�jf`����[vP�O�>����S�@g�ⷉ�Z��T.�P��A̝Yf�&���k���f�Y2N���X�����}SJ/��%
���i�8��W��t��oQ�� �S)�'�bw�нi-l]2�8�&F5�DsYg^�MӐOV��|"�>	�+�nO�� ���3��l9��粨�ȓ�w:��w����,--HMs��KL%�����s�e=v����
\P�4�	b�!S�M�#h��m��G/	�p���Yy(4T�Q;�;��J#�Å<Zv.�:h#u����P��=D��*{K�ws N����=M��2�J��`>'dZPw=}H0uY��!��X�,8g�QW�h�5�!����ur�2�z�Ih���z�O�J����[�����L��q�W����RxCh`�����%֚euj['����Z`���v�щ{�Z}x�%m�ۛ9W�Mf��d��Y�:���"���&�482�#^7HL��/Ec�Uf��h�tA�B�e�e�?{�?�q��fȔ��x0��t�==w՜��EfD��Tn/f�-�r-��-�(O� �.��&���
�R�����z>u�/GNs�����x{M�EO�:��8�I3�Ā���	���uX��q$���+ȩ�a�*�+�h���v��]����1�W|��|�ž�_�ה����i{,?�-OlNljբ�� }1��}[�s���/�� ��{̂�Q]ߙ��yq��o���Vs�=�g8d�u=���έ_��#VX;U8&`�?Yq���}S���6s.e���ʃgf�vuTL�f8vuE�C��<C��|�8�?�zHC�C�(�Xr.e�׹S�N��{�;N�{�	<]õr��e���Ӵा��ē�ȼ�I��Ri~�'\	���w�(�K�?�z_��+�Gr�Q��F44�>��e?�Gjh��&Wjx]{��A�=o�2��l4̥����o兲Z��V�}x�ߺn(�g�Ҹ���ܺp�»m���Y�yƔKUhثOE�B�r
5�tFR-"�>���Z��������x�������B�+�iZÖk�{��T�T��~���[V�`̪�qa*�RM,~����uy�Q�"�N�������^
xRS���e�����Z
�&�Z7b���A�;�C�'��nQ�L
R9�����~�8]W�EC��q΋/l����}�)�5+���y;�/M��+^��%K�T�8����7��uX��i�xQeȻ��|��p���d�,�"�	Ƚ�!
��T�V�^���EAIkjsm�3�]��m4Q��|v�{���{�_�<_^�����>zM?xSz	��U*�����;z�T'C�{��zL��r�TI�,�a6�S�&�_k�5<\Gƚ�Y�/A�w`����������⾟Y�ۇz)�3u����?��U8��k��1��q-�K�oI��p����L!��V`�1�|�������d�Jׯ���ʀZ�Z�8.�*4v�z��B���Sz�b[&�����'�YJ�w1�	�G���,of��$Z�Wb� ��n�,.��֞#o��㵊�� $� <��>k�����P������ah��1�e��ۯR���1-��]O �{8�<!Ǫq��+zˇ��V�(�=U�JbZ��ԸZ���mp�ڋ�5�%= �xn����*�$���k���7݇\HQW�;v����ۦԐB�6����iűq�,���^�i�5�`ԯ{QqTIu�cw*����]��@�#�� �z�H+�4#m(E�aX�Js�6��(c�0u�� ���hd3'u���<ت�M\����d?�&�?���_�+�6�m���K�iF��P��	��bL�'�����3W�̗�b����~�`�>K�w���B�>pf	�ˬ0�aGD�\~�A�L��WR����yR9<l��?����l��(
��reS������l.���42�:�i��Ne�/H��zi�HM�C�pd �K�Yٝ�����:��1'��.�Ut�{��	���M��l���}��0�{�R{mg˪(�B�����R�֓�B]�u61��z�=:��S�����}�n�D� #��[�ǩ+���;FY��8��]6���L��
�9w�M�Qg���D0C@C�]��h��y��Q�᥂�r����<c<�ڐ�ܑ�+�ێc��Ym^]�M���C�g�0@]oz��R��o[U����[x5FL'��/�Z���Q0�+g�4��4��8�|�F<2�!��C�u�I�E�<H����Ť��u�G�g����H���A����ь���=��?���gQB��.�"�%	�#���vA��Q3�'UM׎���u��N�MՖp<�s V�b��pV�ƻY�7>��	�,2ŨљH���e�����$Qn���7�#�1e�����vլ�UΥ�좭3�bM�U����Tj��ߟvl"*�̓�N���@q�bפ�_�������{�V�:�u*� M0�*�)�G�����@�v���Q����b8.)��ݘi�Y�?�˃�Sr,�m��J�5��F C�����6��Z����5��R�H��|�x��o��= �dդr�c0��}�ʜ�$B{N�!�Q�Cd������2r:�ڠ�%�G{ʔ�2@p�?��P��s��"3��}�G��Lw�l'���:�gKx��.fȍν�14(ʃ�!��B�.��ʻ�y�����~�F�ZU�n�fj��6���U�����Y�M ��@���+�68�e��bQ��\�m�S�h9\J�z��y��Qx�������WM9��$h�^9��z^�j%�k]/�-5"���Јy��J���3��0���lO�b�F3_nt���������w�o�2\-����5�H��2[��&�"���!�ȁ>�4�b��pmuHH}�źW"��X�iU�N�����,�$���e��TkZG�o����ը��Ö��ٮ#�rFû֧�U,�P������6���xhQ��ѕ~+�2�_f+*Ɠ�~��L��	˺|Y��u���y�]$�]��)�75���V	�dm�c��߄�w����!\�|�v <�|�U[���!���x�h�>�s��/`b�&&�OD��L~�!��g�[���1����J�eͤs�?�pl���N�i9.V���/�*^w�:L!r�DUL,foDK�-籚7�����e�ۨ�\�7�& }��3p�9�8|ipzUg�S��p����k���[�7�xSh}藃J}�S��s\R-x'��Χ��W��xH-4pX'":@rVo��?�ʞ��V%�]l��feI��7�;ўbP�;��#ʠ�/S)\��c�6�$.�v-��Ŗy(����M0��a������?���>b%E*�I�B~�4k�����]�j�K�0�	Z�L��ai���Q�,C`z�x%.����\ͅ�"�i	+�~st��O~���$!�0�\���P^4#|� �Q���>���3)%����N툠'�S1��@�bw^��=?�%�w=�ZN�\�Isz��V�;����Qk�c���q���T�=J`(��n{�����H�a��q��JE���i:XH���DzQ����)��Xy��9��h)�uN��[[��i6L�s�WѦ>uL�yɵ�VG+dB���"��3�
Փ�2��`�ݝp�z�;���j@��C���%\M�Wj?��~	onz���Ye�p���w�pAi�R�:���X���f?Q�M`����0��<�
B����R��yTK���]ZV&�ӕ��"Ԁh�"��Y�@�w���#D;�e��I�Z�R�oW���4�h:��B�5�p�$IL���V4Ũ$���Ȕx�@�U���ԋ�_�����O)�1����e�d��`?���e�눜O�c��L�C��@"(�䛆ⲉW�~ÀM�ܱ+�{��`��Y���m��Ƀ㙢Z�r�"қ{�L����G��Ze󰤁?�y�ev ��XT��k'ND�v��%g+�s�o �ݣ+��n��i��� ��԰���K�M��o(�(�Y��N�����b���Vmh~6�bi�}<'���c	�Y��5
�d����墄�����!Cr��M������0����6Xc.
�bK�������u��.��A�AA�ܖ�$���7�[�N;U�B�丘8�Wr�,�h�iX&�n�e�D`��~���S+�*��D�0td�h������6�Q���?B�Հ�6���x\��)j�;BX��&���@���%�k�u�J��"���o6|��P��5���E�O���B�s7�" ~�IL��v�y�v��L��I�;��iG���[Of��ѐ�5u��HՂ@^<���<u�$��� ��Fqv2��k���e�n�ΐ�L
�\!������N�:����:�~�F?�M'2^��9���w7�Ь����Abj���,�6�7�B7zŇ�~4�f+fsx�|\�W�/4�c��?2t|$���Qx��h0R����+,�'�x	.p�� ֈ�޶}��\3uT�Kk}�Ӆ�L�
)I����۟k�D��4? �-��!��؈�p���4Jq�lb�v�c�v�v��ת�N4���9���{rw�U�5ޒu\Mt��k+
��������M�Df�$���f����Vԯl.�8��i\�W]�$kJnFy9-sQ&������Ep�� ��jw�7��m�ڷ��P�\'%�{ʩ�D	�@1B�
��!�Z�T�����o9�y9J>#��b+0��	|`'?�ڀ�G�\�茭l� ��褊��(轑�"Я's���Y���r��/i�A��Ѥ�&Rf�B��~�I�g�N��`�@�D��6Қ:3UN�	�j�XEC���V�5��>ۤ��]��']ltv�B���ʌ�H��t����(8�d�~�6��1�����k��;9Q��\X~�� ���¾�B����Jn��ǋ'�w�j[V��s�RG#b�z���A��u	�7"j�"&;���A�Q�j��\�������pDR��?|֙�.�$���0s�uu(�*1�.ܞ��l0�pZ���=�V`��\��}�V�⅝�k�/���M)	�ݯ����vgq�HMI�'�8h��%���a�-����k񸁺�-v'�uI�����r��o �\��OV7�P4��	C���U�H@����s��E&�H�?���ǲ�S��a3�:!�tw��Y��@d���[�3&a�Ѧ���-��[��G����z7!�5�����Nu�[0i�\���-bo(77\_D���h��N�wNnd{����y	s��t��eR�����/�]k�=F���&C����n��(��;pw$���xY"�M�(�)�> ����$��ՃЭ�r����0����_�#p�0��Ԝ���v��0�d5g�;j$Ǐ�����S�nA���
��Q��8uI���҃�Z�PIE�Y.��+��s(���B���
��8u�Ec]���4ut�w�,�M��1�\�(���3��������������1��6����i?�3���[|�i�+o[ �z�tmfḆ�w�����u���4�K[�����
%�nm%p���\���ZL��#�ބ�ß�^j�����18�	)�l�I<S����̙�Ǧ���b �]�1�O;5 @8�5�?���P���%�&�l�X�#�����H� �I�=��F�介��A�,�k�������x�D�iX���-��1Ã���l������B���!(�[۽�A�L��}Ș|L�{�G�7�|�X���"�#�z�=�`u�[����6n��ˣ���ΑCg�)ΈB�М��(r�d5�6�3?��)VW��D�
ɐ��D��w����G$�1t��X3���w%�_���CڕƗI-��B)ƞx��Qˆ���E���ÿ��c9iyHJ�w�D�c�Zs��'D0R�IHzK�܊oD�,(;�i�m`[4]�-`$��֛F�����������s����i���ѿnJd�z߈6Q}�M�ӹ'Xd�)`�=����Tv$\v;IA�그\	�zE�z@<��Ӟ�v0D�#&r��＠b;�j�qGo� �$�Ūr����3�b���G��Q��@�VY��p�^�ت���8�<P���Ͻ�� B5��pb���W}�GW���q��e���\T<M�V���z�y�P�� 0kK���t�4|���D��b=?�
Ǎ��ʫ�ڥιw� Ԥ�oߎ"_R�ɝP�k勚�CJ8� �v�5W�&�qL�4�ؙ�Af1GA;���6.~�j�2DRŸ��m�b�,�U�� K>�d<�g�L;DH���F��ի����J�����9���}���-uE��"?}�>|A��OK��n�aYX���/��������gc��`�\�+�\��!C��C=���v�e֔\�c=x5���y�/^�DC��N��K���A�$�q4�V%�az�İ)���-�K�/��7N�:M�����W8�#�=��KVf�����\����{q���%�`��!�*��q�����V�����oN�L
;ی���r+>�F��[�;����7F#pZ��8\7�s����ĉeI��4�c�0�K�@yK�Dm�Q�[���)�������eFT�s=RƜ�p=Fߩ��OK��
�Ɩ�ā�7y�J .teSGR��[T�_�BU��S7����29�.���a��QLf"D��'��f��gL��>�.r2�L$͗�IuG��nV&d�/�셯�:�À�{����?H]#������v����޸B=jX@�Z��"���j�N�М�b�[���.x�E�P��n��<v���>��s��yPj`l&o��X�tU��|�M�̈́B�Ȏ`Z��F�a�z���z�
T��9t��l�Z�A�?�rN{��u���d�0$���h�G�6�vzGaV&9X�=�נ���)%�B)vhZ�H'Bm��	ߐd{�M�z��1�k+�/��]�B&���8/��08�6����(X��vWDq��J�5��W�����s�L�k�V���M�]戴E$�{����<(��]8��vy���}��Z��|�;Sas�I�wz�w��X[t�BG6	Y	z���W�w9ז��#2��!?���p������s֗��mU�� �` �"r"_���
2Q)X�'��uA]N�.^������PXk��.� p�>'>���&���?�=!c�f�W(��أ^!��h�'�F�a5>0�*ă�xt�>������y8|q@�V���
Ǽ:~7Va�*���t $� N����: �k�� �qJ���t5jB[M&���G{�9�����\o�-6Ogm���Z�q�[W!Y�kuF$B�C??�G�ZC���1�X^��#q�W�u^Pb�_i���K�q�V{'�?��$�\�(?�^+��m�� �.8��ģ#�׺�͑NXK�x�ac����P���S]ʧ�z�A���OQu��@�t�����1;��Lh-���6�w�w?�y��`~:aڅT�j{,�Y���K�پ�P�U��B����J�SV�Aҏ�H-�ǿǒ���t�i����m�)�ҍN�Y^w���X7S���������������ohvR
�q��H;��,��U��'�����/珽= 0�����Y�vIv�QK��}Q{� ��:��}�/ד��ƹ�O�Z	m�#�Oc�Q�J�IM%ŭ6ܙ�͏]�A�����V�6����q:qd�D��R��R�c|�-�#�l��I�������uR��8��>o�e�6Dl�����i�[�J�sl�a��U��i���*���MZ6������N�:	γJL�`�A��i\��L�%x��R�I�!#ڜ�g-:�|/G�9�hY�nR�����P�`A�8[3V��$������bv�7��~欸(��3�9^�_��h%nB0#���'���+�2���t�� ������-"��n�5z/�(}�꤬T�FЬh�Ə밖��s�-WoS��̰\���*�5�����;�0�0�bC�{w��G���Ǵ�3O�������+DG�oP)��'oq?h�]��t@&���}��-�R�����Qt¤��Դ�h���X,������ɉ������fSA<A��ݟ�����n�����C��WU�3��T��0ʽG�&I��̸�A��Oھ5tE/w�$B��3�:~�=e��Pc4Lo�xp�J�dX$B���cy:���?�5���Ы{��-��qb��N����BA}��y}cئZ�պ�Q�`�6(,�CBltH�<b�.�-�<���>���OK�A>�⍮n� ��{=�U#s��#-��k��k��ߵ'4�t�"�iR�.u5�R���<�0c4�l�[fB�M��JL�e}NLA���&&O����F��.:��V����e`*�V��!�n>���j�̰�KX)n��D�Sd%�`��GD/ر0�.�ɫ���z$����X�]�\-�X�w7�ۧaJ�g���n_.A�E٩^��L�p��T,Z�$Q�#���?�kw�/���3Q�gP�̠��r��-Pl�{�������/z�<���Li�pa\1��I}���os]F���9�w��hJC׋���C8 ۬\��dj�8�,O?M9$��Oe�W�Hy��1�ʆ6>m�b2��=�f0yT�]�R���Hy�ח}��1�9r���R�{#)h(��@՞Y��m�_�ޝQ�j�p��p���<��e?k�j��d	��^1�`�m��ݒ5R���H���ݵMOb�)��w2���ؘѕA���?�c/(��V�v?\xF���kWv���M�1?*!2��^��8y�d�3�Xvȥ��v(��+h-�md��La��2xq.�	��� (10Bn�&�>b�o8�6�06�t�޺���3qg��D �5t��J
$5�hQ���c [�f䧶!r"�J#!wN�	���o[k�����;/���(T����˦���?Ħ�1�x�	ٝ��O�]����+�( c�#�{��'��}ƨ�%_�Q���{�����VB�z5�4ȓޡ)�=N�ks��������j�L�Cs
əP��9��'��o�#�U��� I�k�M�MJ��.gR��^Ӣ���D��� ��UD&֜�/��Q����'�{�vYv��E~���,ewԆ���i�
���NP���O�dk�'ĭ��B[��=�b��U@+h?B:�>���S��>s�}c�7^���Θ��#*8�vA@zM�.��]��p�_ ^tr�o�R���{՚_���	�6�<)���c����Z-��bP$-a��l���h#7 ��� ���V�f|�����qٔ|K�n�d��7�w������:��~�kd�3m�t�<2AJ�������Lb�,�v���b��sE�x�i�̸,F�"-�up[2(�]G� ����^\�+a�NK�� G�/����u#�a�{��A~q߸~Q��Kx\^&�r���O���wm<d9Ƒ�qNr���A�晇Ӳ9��¤���R�,#d)�IPW9���[������+��W�t��d��l�7�a��5#W�j��(��V�ʬC�d��ZL���*a|��w��
�%`^���Gp�0����ߩQB K�Iѵ��~i82TІ	��o1��O�x/�U`��5vs���O��% +t���O$��f�]��9�_ .|L�<�ZX}�r�֬�|z�l(������E�ʘH��[����Í��}
�^�؄�"��)��Պ���281{�C��E�(�i�0�(Z@:���HQ(D�ؘds��<t]���3]��Qc���"RI �v��r�Y��2�'~^[o=V���Kae�_6�/sS���*�Q)0�'g�� �c�c��_�C����L���-����8�/@��j�!�as��k�#���{��V:�K_z�<$��!W���pVK�<��,�b8���>��G_�8���=��!`I� lԛ@�ay�Ug�c��G���="��i��Gɹ;�ݴ�XR3��n����`�=���+1r��O0�"��ɦ�>݉
�NJ	�7�n(��Q;�2aް��u�G��]��W���[�m ٿ�i�/
f@�I 0��h��F���f�����
�.uG��|��;����f&����t�b��/?C�U���|y�l�������eI-�\2�F��q��霥�PE���m�#¦�M��� �J�W��N�������R*qi�Tx�c�k ��y5�����v���X�S�I�-�pqV�s(N�ȴ�	�6r��d�wÄ�L,t_�ո��L�<�ə%>�L���l�p�7�{'��QZm�7�]N[���j��Ucl�^�۬����m�c;�z�OD��"�rYgl����^�)G� ����u2�j��{z��ei
'Yc����k��D�&}��üJ�?�1%�D�?@��)�sW����7k���P��5#��H�V����|�"��^m���-���C��_�����R��#j�XU񁩂������n�n�W�z�)aJɴ��ǫ�{9~�P�\�+ˣ����(�.�< �$d?���e�
�f�h��Y�|#A��$�o|a�Y��:nQdn���.�'NW��$����LM�6!�3�t#	���;
��·ɾ��hkѫn����s�z�w�l�k&%S��������~���
+6���m�����d�Bh5���Q	(y�z�5[T�ԞčB�R����
{Nu��Z��*���%���{-��t_>8ĝ}� �z���1�[����C9�<+�D+1�iJN�<�_t�ʐ+9�ӽHk��wIb8Wh�:�:�;��	lwMXU>�m<�?�S#���)
a�l>ڡ-gH�@m��~JGV�W7$e>�LZ��e(����"͘�'(`�R�#�1�!:=� �޹vДb�_�#�/wҴ�(j?�H��~I��Pw�S��{q����SmL=���P<�­rRY�5_��4�n��BN��}ʮ3���.,���Ns4�N\�&P�FD���'W�d��J��?��g�,b6�WQL�ر�����Dt0n�c{P�]IKOBG�S�l�PW��I��Xy���Zx������!5u��Q.[XX��o���7���8��%�q�1Qu��ϋg+f���;��u�O�[P*�Z�[�m99NC�g��Jy�2��w<�e0��D�R=(��_���	{�<�����D���q��8�
�}�����!WB2Zu[�pk9}��� c�w����0Yf��}��蟝L�$.�=^D&˯�b�c!*"2"�8x}��
��a�9A����+�2w"���O���.CD��BJ*�A}��B7�:R�'_����b ��kı�!C]'X�&�uVC�?��oj�H6=ٍ5y�)�}P=����fJi����
?�UPdP,˚76�h�J`h �kF��hw�����lh��s��Ќ �q{ɭ�2���}�DJkV���`d��Ȇ�K_F|(�љEy��:i#,n�"�tѩd`�h��\�����7.��=2� m��6�}ğZ��G�{�K*������#v�^��OS�Z��:���<�'4A{����a��2�r��qf�2��I_�����T�)�{��.uq?W�%�BX-p��4�j�yRx�Dq��eW�ˁ�rdr5Ma�����,~C�����0x��[9`�TwV����e�E�D����w���eA��!�r�u�a� Gpm:�ޫ1A��G��S�q��<L�Ͳam�N��4S.Qs�SKkW{��|s�`��:��o�d��Rʽ�u�کVcm����b��w�Hᣑ�A Y�Ipv�o�S��7wl�'��M���i�}�P�������P�x�`�f��t�ʯG�.���T��Fg3^�����q^ֻ��>9�jr�Ґ��W!zXBs��'Si���˺��xR#tr��*��-觍�vY��(mN89o���s��lk�<p䌖;6H�K-���"�)e2~*<�t����	�?�a_�Fo�A����L���M��Fk�h��p�=x�BK�2o0LףC	��\r���hCv��C^��Txvx�KHw�nu�_�׊��=S� Fi�zp�K�`]�7_�_	�u�b5��
��^�l�9[Y#l��KDJM�E;�)e��H]B������ S�Ixm�yU�q�'*L��|E�j(���y�_���i;����j�����/m�2x[:w�ٔ�Z��M��SW�UC��<��Z��o�rM]����g�O�CLOϴ�y/u{�q���(���LBpA@���؆����-Y_������褨B�]|W�OHEjN�΂҄�y��À���p*Q������S���|�1�عy��!�Mj���TX�L�ɗ��������e&T.���؅s�����1��'���kpӁ�I�}-|q�U/φ2�����{]�*�|���,\	:�T{sMi����E���T�2�C��~�6�w>����ţ?DZJ�=w�L���2��'�t�8(AI�?��"J:v啝�4�����E�~�u���,���A�r��F�4���0��C��fπ<?_R�y�Pr,��3�_�
���S�v����:������^�m�%h���M�J����ѿ�G�e�";5��%��Ɩ�x�
S{gQ�k8H� *����O�����8ME� ��m���5ldJ���c��5Q?����ߝ�9��4�$��,Y�\lQ�44��K��?J����g���/]�-:��ob>Z�[.<PPxO;#���'\SԴ��F�A��$H3@��1����fJd��04����魩B=�9�\V!1�$�> !�����W!�7�0y�b���n��}���>�>���;|�����:2Ug`u���R\�)��	��i�v��\ȉ�Th?
�_�M�����N�Є���X��Z0c~S����%	QВ���Y��m�X�)��羿��Z���9�mA�l�d�a���F=�Fw �lH��u����)���.?� %[w_�Ⓧ�1:���C��u����]��g���{�YagW�{ІD��J��X��{�ï!\�*i �h�P�F;�U�#��>/�V��i�F4"�76�����lL���diXO��:RâyL*��3�l+� �?��ޔF^D0�s�
��+t��_��n�E줿bE*l��Q+",Q#�g�b��Lv;��t��W��Y~�~B� B���2����^�6i/�\6V����x��H��/�ag&~�pI�N����`��C�D�����8��17D����݅�����[�����~��#�X)�]�^y��3JB�&���n�erU�95?���*>-x;�~|�Х�ECD�^�'J-��YI���ƀ�k^�:1�u5�F����l�Fb=X����^�#�9b�����D7�Emj��nw��5��ۯ�E�o���M���LQ�N:8^ ��7���v������5�76z�	�eD�e4M7��v4��3�����=���M1)ę���}�����h��vˤ�m�N��5���҇b�!��\���|&�x��ք���rx����Z�Mi'�����-6�(���6tKд�4�9 �{���om���,oA[���q_�wK��*�ʼ�qn�.ũ��B1s�6�X�$�諭�5(���YM�)�JN�͂�؊7m�m����}��G��ׁ��!s��_��6�O&�'*����s��'���t#���QR�1W������D{ջ�'.�l��>�@�P��-L�L������)��U����cn� ��lm8��UX�},%v8b_�)q�#мS����P��jѷE�`--�r9 �Z�6+�BA��ל�Z@ts�������w+��N͚m~"���4����QATj�g� �)�������靓3��|į�ȁ��������[��t仜�V���e$�y���ŷ�5�i���y�q�����)g-@o]=��x_FOk������4�=�K��U����<O��@���o ����U��K��~��.�~��h�7�]��ܥe*��_�wU�W~�O �]������[ &�g���4�c6� A�u(9����>�C5J�mw��DwǙL���wi�`�� C����X>�>=2u�'�k�g�haXg/��x�{�y����h��Vz���;/Уwbk���#��x`���1n���(��)�����,;�=2͸�ǜ�.���+z}a�+?�Y-I�Y�0@�i(D�=��d*��ˊ�1 ��,�U��+-@�@��Wu���.���Ӳ�#4�����K���� �H)�王GV�_"�1��Mc����`@�����0`R8)r0���ug�M��<Us�Fa~���ԣ�زl�5U�b�a;��$9�T6=�E��Ju���$�p��8�ɷ�nJC�*xs�у�H�y��@���y��?����^��}�2
Λ DaӬ%��3��j5�����͔���i:l7����Cw�1��_(d5�17���;%��!z0�j:���Y�[q�%ܻwiV�ʚ���n�E�V������:)(�S7C��1��p�~Wpm�����?_�����r s��g1�?�+͌��:A� P|�
(��Jj���nLB �2٥{jRz��r��Y
�<��������t,|A�K�Ь�]�T��_M�Bi�t�.Y���ߠ1'��Ѻ��ے�:R����2kT�!�G�,����޺4|#����> ���~�f��d��O�5u|�(��0�ƨ�
~�dԝ	��X7��)��K�ݻ�Q>��1H�-�65�*JC5�����4>/�$3��f0�9a����Cn�.�������ղ�*E�z\�[���i����brϼz��T�ܱ��2�����.�� 9Db�
�A��uǹM���1��Q4X�$��CLڄ:& .զ��Vk�~�c�<���P��t���; ~�a��E��k��_&w|]�6D�U� 3=�f�m��q��.�/�vU-�㾽��Ulg/-���zh��8�z�q��qHx#+��$�a��t��A���\�{�v1�aޟ�]+�S������+���O�I�F��^h^/v"����~1���c�#D�}���Jj2� �
)��[i�⓽i$TG������E��/��a*��M���s�猵mȗ�5��9v���H_���jl�@�����^Y�7��!Y��կ�����z�z�)E�C!��|��{ND����9?��$����|������ճC_-���aT����a�y���W5��vv;�~H �#�.L�]��(�H͝���MB�^��t�*�P��pwuW�@�ۜ)�A��}p�� .�n�1��&��j�:]'�ޢ��1��M`�������g!58Ї~���t�_���	���Z�-S��B�T�><X9! �S)��i$