��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cЌE���MuW�H��I�Qʀ�v7���4p_�����Z(���ɠ��h�Q��x��x+��lӖSU�ؘ����R4���Gl�?��Xٺ)��"_;���f"���d��/�Dj=P6�z9׫}0�Ln��R�x�p�/w�bkS����.�[�D����V}�X >ɛ'!=wٓ4���	�X��h��t\��Cj��~����(I�o����d.]�0�=Ts�u��Q��{�(��>l � �A�m�A���'���,L0��E�R��R��}���`���I4$	��+�Y�Lp�D�È�
ߗ������\��Uֳ=nrqq��Vv�D݁3�"�WA9��;S�Fj]�� ���)�~������=���;_B:������\�9a�Jg�E����v�텇tj#��w� ���;����E�ϩ�_� ���i�DZ~zNy�h���6@h�2K��	گ ��66?'�L&�6�b����dv�z4��sQn0P��r?SVz���X̳w%��ᱨ��Y�H�Z+�K�z=��M9�<�g-j���_�������b�%���ߢZ͖������;�)�]q�zi@������N�;���A
C�N̩)�H�<h60Oq�1�T�a49�<�����>��� +���-^�J`w�t��mᕳ�6�8mOpڏ�8�MJU�^�%pOf�kg���� �t��ߎ�5�3j���h��$�M��!p���77��%�Qb��F�P# ��A\���P	���ڶ��W$�h�@z/��G*V��n0K�L�pu](�!��}���a���T�G�3�j]��-��e�!^b?�}���ė�h��D�T*4{���z)��3��

����κ�1sR���nH>� +������"��-g��(�L���47Qa�,)��)�>8w{ކy_u2,��&��A��s
���>!�Iթ1���{���Џ.-h1�����kPI�
�b���My����,n5ꑳ;�a]ҁ_�u�Dl3$��oQa���lH��x�� �U;j�&{^���/�|�������ꇮ=*��6��
��TX�z1t��[��먙�N���9���6�_�'0���gh���6�+٢
���,7��M�SG>��1��q��J�0�lt-�/�7���υ�gZ���MW�i����Q��[�~�.͝�'�>�&�Օ�[��!�d|yס@�=��GT\� hO�lW�7*eK���4環S|�U������#�$�~^*��/F+I�+����=l�LR�&����!��ܭ��3qh%��iS�<���m���4#Dp���ֵ��0�" e5��;�N�jA��ƀ���T+T1Wc2!+|��������c��s�O�1��I��_�=�jN��%���a{x�+��}��2w�����*7_��G<��.�:×�f�is��.GF��'��3��6)��\��l� 2��P��i4KT��\b�OՅ[鞔�r�7E�屧�
�LNѾ/K l�]���*~$�����S�j��Ml<�2�w��̧Cmn���p"�q���O�\Q�^'�$���Q��!�3����5pͰ�c5w�VءDzkC�R<�}��.���cX��tQ�[v� ��W+`yiŜ����ER?2ҳ�����x'|��꺄$�>������ʊZQ�}*�:@%�;;{=ޟ_� ���\Q�ê.vđS����*=�_)ن�m���h�Qӌ�j�8A�O?NY&�O54=j��<a_���
��=i�� n��i�6�L%�s�X��v.`�^�|�v�l3�9��2}�Bo�E#j�K�7t|⪀�$�!���6(*1�pψ���|L��Qg+�hqM�k�s�N���?�cCӋǥ�����#	� �E�)�&Efp.Z`#N�'�á��E{x6��ʨ�]�jb���!����ї��� ?˜�-��6F���)lk>��5��0��|+�mu�v.[�?x$f8�DP]-[8��ɜ��=���M�R��^n�wĖ��=/���H��u�#1��1�U���_~W��)#��n"��Oe���hJo��j���� t���{BjH�n�\�l3�U��ls٭������3���F`WƎZ���x�2Y�C@ �>�`r+�2��M�53��'��O#H}Z��և!�U��Em����8�:���g��p�ݖ�*�IT�m�|ztT�8ŵ�ꟊw����=��:( IMQ�.�H7Tw�Z�;��������0������ߠb�r��FY�	JA<C��:��N�vҌ�6�4# �.����Z��ܸ1�*�w����~7<d�X��,�<��Xe-�水9-S����y�/�;��J�����n���yGrT���j���<��"n��LO��,�����	�j��iោ)��_Ir�lĽ��*���"j�:#��{<��o�buδW���#�N���wh�às!���T�!�8���lҾ�+Q�{z�z�<��2D�*�?���q�Q�e��O �ʙ�k,�eD5�/J�	|�Q�Σp3�2�(JT�~M$�t?%;�ٱ��M�j+�fDU3�
=���n�*�kz����@��>���F��P��Pg�shZ��IZ�ط-��/��<yoHZj"P+����'���7���{����.�q�O�}��y��@y�¼�:�\t-@�vDF�w���d�`-��K�)��?i}�U�	]�Z��6�F+��9��Pf�Qa@��Nz�nK�y�IL����,��A�o^�ci����obFP�96�)���2�xvXP҉22��������J(�7��Q�!t�1(iن�D�%���2<2��� YvA�1���#`.7bB�L;G�(������07���q%DlX��3�r)wH�,x�P��٪s�K�[���HD#�ޚѐO�5�֖
L���\��4o�ͽ���c=-��~��
\��V͋dz��������G`%G�|>A�fp�m1�Ԅ};��H��\�H�@
�d;�-W��MM���N��" �q�mm����?6���ݹ� ��p�9]J��JTӇ���2�X�k�3N�K��¯�6G�H��]��=xc�w��|�̍�,Aa	�i�8�>��2�}O���WV���q"��XH�m���ǶAq��ѧ�?YqW�&�p�q��]WT��.��x]��-��4 B��s�8���UP.�j�U����9�U<��[�2��J�d̀rpw7}G�|H�Yq�`����
N�
Z�^���SȔ���-���B�5K%Z�b��wuu��.�9�FKp��5(Xi�)�g�����HL`n��CfB���|����m�X����K^F��x7��:bD��/�$���ZiǕc\R��vH%����S���@�
F���k,���J?��և3�_��ͪY/ɟ�~Z�0 ��1<�dPD�<*��9���c�� ���ф�0�%��K.�&�6�v���i��.Q���0�I Ax� ��F�g������4۵7���S�K�: Z���U�(�,#}�][Ѳf��:����`������u��+���{��P����D�
� �*��&�t.R�����@M]�c<�K�P��%��Ud_�M*��菞ڣS���c���z��(��b>A�U/+�vO<!Կ_"+r��	�4�����05��ao��s=�G*�V��7��
C�	���<噉%�f$���4�qN�rI^L��̳~s��J�q��!�D���F|tc�b�u�C��ɩ��.����B�,�#[]�8���t��{q��l�;
c����hj ���⮍y�s�{%�Fr9���A�3~����"�o3VNQ�ԀT����`�Lq7T�Pw�/E��Þ�Q�RYV&���OY�&"�.��E��l$%~�=��6؟c�!�ݒ1Wh�&6ʔ�$��Vf�40w)rR�p�ɖ#�x�A۽�޵���xK� ��Wfrj���ևY��C�qz�q?� �m��h'��v�y�sE�qzvs�[3}f��'�|W$5�0^�jx��B�����O�Q���x��+"Pj��^*���ɥ>�w��F< |���B��DW�� ���?�\���n��&S�X[��R�sϪ+qY:�!?��?��^��!E]�{��ZW�=�-��eof�e�I4�-+_��U�Ɵ_�"�Hۍ�0�@)f�������8��3����H�QaF	a��>�d$y���W�Oک~��{�;14���!��d⢛E��WFߪ�<&�_7�q��r����/�V��]XgM�
Z|O Y�2���˪;�pED�6�>/�[Jf�d>)��'�JШ��VG��l\� J@�Ԕ���9ӟ��ߡ#1t�C�P�wdG·HP�z��ԡ�l��j]�[X&���o���R���i��4�-��UN�<����n��2u�r9%?H�ֲ��xMg���K-�����.k)?I�d��q��')��Mi���M��Oi.t�+�k�x�:�k�8��QJ�ݝ�޿j�";�Aa�=u�}V�M�� ���8�������r�QVi4�����>�Ӕ%�n�}���]�Gj�����MHp*���+e����2�����.��0��^�<y��m������Po��Gr"��c<�6B��0mzq'ǀ5#tz��	��="S�KXV�t�.��h��Yn�\U�W4�+	��ܧe�jiŤR6��r�:O��5٬
�H5%*��C�/���X���D��2�Y��u�<3T)������������IƑ'���C�޻$>�B�,Pzf�|ֽ�W��>{��/U¨ �h��SQ�V�4<j�ЬHt$����i��Xl�!/�q9���x �遑ҡD�mV:�-��,S�8u*m0��4�9��QnW�]S���O�~�P�礳W>bX�g��c_�᫏$�F����'X��4v:n��iWfvF��w�aV�����~��(�-=)ۄ��S˥�P��.�:�J��������&K}�F�`�!a�n����娧�{A��4(s�1�lz|���s��⅏n�V�6����+�� /�@Oto����	���;�0�2����m�7I�l�M�>��о�������D����4�q!w��I��aW�����J��q@�����`�����vf�)�갰��7�>k	s|O�,���Y�d�����z<ȄӍ\N���Y l�R��dwR`�e�? ̎!^�R��1hP����z-�����n�D�y+#>��v�*S�u�\��?�5�"��ٵm@N�K4g]�*����C8P�6ɳ��7�ri�>6F�ܐA�>
s:hz�o��Yהp�2b`�Le����Ҷ�^�TCs�V|ydR�㻪ޙxN�n}���iN4��3�c����Ք6���W��W*�)z�j��֑p�?���vw�b�RZ&=:��X������(�-�֎��W�}<7؞��6�g�v�8zQڳ��{�gC}l���R��L<ޓ��^9�j�����O8ӷ_{V����[���z)q��������4�\r5�8+М�M�o7,���6��8(vA��Q�Y��GS+ZUh�)�T�7��ާ~}�ߍիᏗ.WDR<��%:�Z��	��؈o���(ҫ�?�YҘ�D*%$��Ce�+�f���|�����&�I�pٲ�"ǑR1�����4^��͔#�/�か���O[G*��:�z�u$����l�F8�V��>{����OpP˗=��7�'	]�P!y<��W��,�=Pp�?��%�=�2s���jG�i�r͊��X/���=A��FM֝t�H�.r�|���\9�rh�{2��JF��Q�EfR�M;\��������ԏ�q1�c=�]����{��q�`��;�i��-��މ�ݟ ��sD�ƾ��u�0L�ɉ,'ݿY|M��V�ć�lTk�؁�����K_�pp��:���z��ɮ2���^����[��в�R�4m�������M����\f�ayDQKw�����gf`��a7�!i*[�����3l9ku����7ݏ�61���� Z���D�=��Q�D$�P�YЍ��p�H�N�p��N�(5������;.�-f�����,���w�ndN�h$>4A�=�y�\���;�,�<�,0�Y�[��&2=��l�����{ؼgK��	G����0U�V�fg`+�^�p��ؓ1�R�S�����?�~�n�y������'������P#Ѕߪ�pE��MDn��SΦR���߼��U������=�A���gy�Ie���{�W�e�	3OY�I����
�����,�.�
c������l�w�L�7��j3�̟��z�Y<�l����P�S_�D[@'����ђ�A���*8]˞�$]�Do�
0��ߛ6<st�V�@����^��K|0�),��!0:G6ٟ�P;�� �\�^�D܃Vt	Ѳ�WU>VIdFQ�P!�v��EZ�ƅ�4����#��J�&k\�Z͑尵"�!��鍇+�7Pൕkޕ3��g��rx�5��B�74�Mf<Z4��C:t%��?�mY��4��J��P,'�^r�?� !����H-��5�8x̺���9-�F�C���nv���|���vU��2΁F�v��!�^w¯��z������P�Aދc>��{]=�{���\,���2JLne��Ēa��0�Q��3V�0����\5�S�A���V 	��</j ���C��NGR5bV�쉣�g��)�������i�K��C0/�"L��@��Ղ��B8/I�UR�~��(B8 �5��}�(���8��q���ݏ?sz+g9���R���i�\����E0b8d����2:�D�qn�s%���fiYU����=�:ͨ�w��wh{�h���8��w1���g��$���WM�A$E��F%ZT�����M�^\|?�z�S����6N���#=�t�
�$73��씈{���KjX��_��6���4;ӛ�����'����kn?F�D�^�Jg2��1�ȩN�轷-������ʺ�5$�@7���}�!wխ�����瀪����T�{<B]un{؝w*���O!��ٟ}]]�8���gQ$�*\>係c��gn!�i���7��Jk�4�B(E��5�f����-��Gt���&���(�(F,}@�/�r����|�rQ�"ג�Kh��������4�de�\ſ�$(m��$H�FHR����?F��"_��tBw�#�J��Jj,�<e���'1TA��h6����������ö�*�%>��3��m���8�a���	��.���8SDE�~���>�ꏩY��Y3D�6������x=yhWB��
�ʀ����ᆾ0���sQ��i�'n�_N�1{i��̆<�O&8��6�f��~��漅��v��xb��1��(,�no�P�֢˜�ʅ>���_�"�M���m��!�L�A�4y���ʢ����s�M�X;���Tm�$���J��q�����7��A]�w8�&�N\�=��F�����p�)���qvf��ݰ?�5 �2��n���]���cm�O*��e�b,�u���="�,��dXx�~�^v/�f:��J�j�~�ݚ��۱�Ču�B!��u�oP���F�q����e-��q뵦��av�-H/\$�cܠ���7��}���
_)�x^��I:���Ows�����L�����C��)��hrR��Ǆ�00��5��<� 6M�:�X��c�k<���6g����.+ld�B1����u��{lD'SWf�=�A]��&<�H�!�F����v�;��$�O��:l�����"/ۢ��U��c�J�Js�ƣ�M��@��?�'H���i���I+�C�ɞsv�J��.�.^qc�����_�!ު�j��m�e7�h&EZ�|s��''D��N@6U\㳙����VXf\D� 3�3��~eY��t��W<֊C�j5UP�鶠��Z�%����v��3��n�� �V �;�P27~��O�4��$�h�H��q�Մ
+��o[�5�2�>��_�Q��<�>�o�4�������9|��K���i�eȜ��MC��BXka��z�)S��T��(����y�����P���:U7�/�����S�HL�f�j�^O��M���u���o:���g�s�U�ѻ�VI &�dá����հє��QT;�lt�(5�ӒU-颸�qm��C&��x1*@�T�B��/�$yQ�� ��W�^!S��yPs(��^�e��3֐Z����jY��m��b�0�b�
n/ �����s�G.����\C�9�Nt{�3�IL���3u4���'JA����{�i��"��[���~�Pz�f8�s�h���b���܈���C@5�q�-g�;��T�b��p�KK�'�V�T���	\H�$��A��A'3��	y����U��OQz���%�|������D�j㦢;���8���g�~v`dp�	钣�#�Q�i:��)��1��ݳ���@�؎�E�l�a�m:+�%|gl3+�s���k�F�H�2:f�w�4u��\�Q��=�)�̐D�ޓT+Z�lh_�f mvO�����Q���AK&̊Ec�������:M�O"c��<�-�:	�v3=s�fd�ޒ��2����	�
g�y{<�y�M�3n��JVb&�`���a ��/A}�L�i�fD����)�E�b~�L�L�FQ"�oѴm�Y4V�ce���<ԏhɇl(���ju].��]��	�����:fɡtUI4�w+�H�����DQ�3fYV�̓���tS�۪�"��L�҉3�'u��&�����L�ѥ�9O߀��H�Ϭ�χ92�����ST�*��F:A�c����D�Y�/�ե�LhWwWHK�BT5Ȟ��f�5����X5��'�;	Q�bZ\�O�x�8f�5*�\uBH&8#ęӻ�Ϗ��Mx n��8q2�x]!1P�f<1��T*�y|`�:�����Ͷ�cC�/�0�����Q�V,�8P�m��V�D,�c{�������Dy�.X�p�5�G�O�c��4� b��p�1r�p�y�Q�m�ۧ8�:C�,k�}<�����Әټ�5�}ңxxl�] �փ�^�I��Fyr����a��P�U�b:��r�ә��_{���E�.FfTud�M����rH�����N�.�������o�ѕRſ��vH���أ�)�+�7X"/}"�q�K���u턇�/S$k���9�M�v�lП%L��:Yڴ�ï��Y�3�x��)����h�����*�A�������N�8���L����tu���}lQrNT���F��֖z��'_�O8��AU�zi%�-H.5|�3�-�}�ŝ�&u��cY�����Gh�p�BB�����3��d�G��VsE�٣�'�րc��|p�Z��*�û�A��	�s6n)�.���� ���]wV�>���1ߒ/_m�Ǟ��H�}JQ P	X���������M�D��h��{�7��K�����Rdz�e.8�~K˵��v5���![$��;}�>��u���e�挝����w�B<y�3ڣ������	w6~�H����
&D�<Y̾����+�˦�c�;5��]iUk�gR�{W��$�c��̪��J�x�E�*6GI)	�<v���u= �C��ӄ9�L��%:�������v�d:'�9��x��-�DY`�Tߧ�b!W�;�NSxl��+߅�YR3�|7U^����Xp�"?��-1�R�m�6�3To��κ�;V��8:��k��z",%��W�)�*�$z�C,���5���+�l�s���O�%�dG�V���X1���5S��8c�n�����G�<�K6����:Ѻ,C�b��.�xE�2�KΌIz��d�Y�&���R�l�p�#A	�+S�(�=�=�?@�7_��Pb!"z�%`��-�4��a$�>O�N�����3��dW"]�jcDN�"8*�P�+ 2�lV�#�:c�f�q���:����I71�T�(<ݞ\�Vl���d��b��iv����p(+�B�m��0�@d�)0�&�P|��`���7�Fg��d;�uZn��1�w���5�����A���Wu
j��B�Ȏ[����QX���bfW|b�N�,In$��Ѽ�������%"�IZ��_�ל�cz�:x�h�$�Lۦ���Ë$�t	lND�G{�j�H�fx5m������+r/*��O��ܳ4�c6ze��`����y�I~��`���{H9v��FM��xo�M6�J}r�U����2��%�M,=��XF6B�^��2h<9�?qYW��cى,*v��Q�rSP�(%8)%`QZp@aC�!�� f�Zd�W��4_�xDw|_}���J���O��I�����&:G����xٞ9�:�Hz �(�x�2Æ�F>�ʓ�R`T�K�����X1�w��g͖��j=|���ZJ�/\�X�i�G�T�a��&ب4�A��v�+0��W�L��\�����<��k^F�4'ht�6�T3��cIe2ao�U��dW\.[v�ې�*y�,��N�f*h��>�i��R�GN*{��n�LR_�H��&���1B�"w(�X��S_f`���q�i��\��P����{D�iesW���V�Twv�P������]�#����	"X��C�O�&�~'��a��1c� ���c�,x�����VA�~�#q(���=�|W�J8?k����hib��#f_�֫}�������F I�	j��l���Kx�TH	9�aٗ��ݥ��`��H��������u��Xm�2�_ʣ� �l;��%�Ӕ�XQb#����d׸��Q>�4��e���!,�
1_W=-���+O���G��RV�@��f�zR���cU`1�B}��@Qz���G�g~F@��gfc6UyMW�>����w���n�s�
��r���-b��xS��bf�z?�G�� oFA���t5��dNa���¼בW���9�*�uڐ;GG�hS�=F+�V�Z�����T� դ���,/>h3���:E?������2&��Wl��#|�D�C�$��3Ȳ8�\m� �W���Pb�|+�r�J=@ӌQ�F6��\<(�4���VO�������A�D��n�Q��:!H�yz�Y��x�o�n�*e�ܶ��[�Ɍ�9yy��u��#�_����g���]C��Y`V��w�� DF$f�('<��w�@��19��S�n"��>��ö���3��X��-IV�e�4�ү�E	İ� 	���3�/��;E�̤�Phw��Rl��!މ���JU�&<��p-Q����]�%�I������Ca��aT��-������ԭ�5�x΍?I���=Kš����&y-�{�P!��k��ˠYQ'P�kl��R�4U�Eq��H�Y��7�d&��n�I��\Ur8�Vv�/B�:�L�l^;>e·��m{7?j5���hٔ2�'zf�����"�!������A�8�k�5I*�6p�g�uh)>��S��?BL��M��\��YκP�$�E6��.ɮ2>�)%*�/ؙwNi�^���^Zҳg�����ru�G�JA�� ������x��Bm[���I�\~s*��_�Z���^�v�Gj��/^�qμ�7�O��/l(9�-I��z����c�X�&��Il7�=�p�_�x^"N9�����'��ͫ��ֳjPY��'����>����o���/թ4d	�؊a��?8���8�I� Z��	�`�]�3�i�I�؈���Q�&ҝ!X��`>3 �t�l���/��S����D�,�₧�S�3��s[ �����:�p���D7��i����]R�V{�>�L0��D0;O9A�x��ڑq�}]����e����q�X�bģ�	0�Tc�-�3L��2t�BG��sa�%��I��~��RQpl��v���6�NҒ�n�_Xq^�z۵p\��)}gy��\�$�5�lu��wJGny�2v�hļ�eX6�͌�V�"�r���F��!��p�����[.�����6Ԙ-�L1R/f���Ŵ�&#�V~�TŚ���N�ya�}��T��*C����pw�R�R	pND �{��T`xWV��'X�!V�����ɝ�*G�e�/ ��\x��,��^�*�n�/��/�	ז�I�����(���A��[��٭
qK������,����9�~Ux�R����
��N�'����7,���u)��ϴ�Nr���3��`��
�$�E������U�O�,Ρ���gn;c���á/��C6,�+��N�]�����]���W}�J©�骺��� �������լ��bp��t��6���Qc;{�Z��O�����ٯ8�c-w ׯTr�Qe/hRV~�6���bd�hnMmѪ��W�@�z��c��dj�q�_����N�A�5�A��eO{=gڜP��Ѣ+B������l��A%��R�0@a5�R�[	�k�KUnmL!Qu��FǕdDr�"�m�Y��W��I�֛@��� C�G�JmV�sB���iOwl烈9�<�mnM;�1��Յ����D��,ڥ�����%��{^�<�}����R7J�bz�@�f��;|�L�q2��5�L����b8��6�3������X�#���ů���w�4�-pDg4QZ�'B*�y��pao]������6 .���R"?�z^�5��	]��XLh De�\�!��+5E*}0�kG)w��x�+��8���H7��ŏ���mٲ��t�n��P	l��M���m��#5Ӵz�<�\2v��u�1f�F�=��"t`ȕ�;�>�_U��: �^M�fJe�!c�O��׊��%��0����OK�,���g6�p'?.1'�=8Y] ܧs����� ��`�3
�T�=��2�ұ�FRl���� Y�Q�9�uZkP�A�!�����6��[,R�R����#�z��e�.h�H�j�M�c�4,���A��������
�	�b���Ή+匢1L���ŵѧ��@�ᄖ����]��q��V/��3>�:�	Y~��`Z�\�&<���9Ar�m��t�y�Z��r�;ƾ�!��Q2\㼺�u#:��P�+���E��d��|T����Asv9���jθ��,�4� _�υ��]I����PA"���}09ʂv���+|���?L��g���=t�Y$�ꗑ/���o�F�Y?3'C�Pm-���zy���R�h��|z�Xu��.�g���#���ǳbw�8���/��1��m،o�lLz���y�j�/b�S��YࠇVs�p}�M!�ų�%b�mA�kk$�.|�0�
>�M�J������^����/7�Xg�i1������1������\�sۛ���l�^��e��-\*R�����x�H�++�:�׻�i}u��y���Bp)4�74��~�ˍ��fsQ�$�D^���:(�-IT��^�(�� H�i3�2����-	��يǧ�ZN����:ω���n?I���wW�vF�Q�'�p�X«�cmﳦu�a3�G�:�d��o���NF$9CM��cݪ	�E�2���2�#�$
�d��b��r����|@��K������W���H�-,�h���_[��[��_bTi�S����k�k�v�2�g����ԫ�rhW�gt���cV��y��(������]�<�]ܫ�+fl3b|��ǵ8��D�A}[��J��	�!�����GZ+j�/��P���Ł��(�r�/��b:����� -.t:eY2r�J�·�?0�ҡcT�5��y�O���2\q1��+�z�DB��Ym�>8��oh�h�U�a�>�%j%�e�%��h�G}X�x/�hs�'r�Y�,���R�r�LN2�"g��l���ҍ5��60�'/����-�1�D	��K7�h���9���N���(�c��kǔ�Ox��GS��&�����FN��z:<�c��0L��v�L��&%�.<xD�*JzC6ooڋ��KhW�S��e��E&���E.�����iM@�)�~z�tV8
T�Ù.��T?���ڧ�]Jg�`H���h�{��
����
r_��̞���!-�5ҡ�}��h�藽��ۏl��b����S�}��� b�_��j���H�x��T_{GL�]"���ui�8sK��ٖ�Ւ�W�kw�\k�����c�gک�V�ʻ��J�P}���է�w>�o`�C�h(��t��}��%u^R�Mnuk%�71��y6������Ү�1���(���@K����1��zY���n��e�����E�8TG{�;��Ae������?�QW`�����ƺ��;of�0	rbo�Ҏ'�7���a�y�Ol�*#��na��r���Xޞt���UQ�0#�9SPV-�-�HL���Ǿy����^���Nz�
����
<N�O�zQ���lq�C�m�މ��:�}�~ :�ف��A���6�A�ՑIh����݂B	
י$;L���T7�LV^cm֦�e�q��;����E��*��ߴUv벥$Y`���nH�EI�wU�f�)-�)c���6I̎�JS�H��K�2�v}�?W��M�f���{��ׅe�l�uf�,1Kk"�贈�i땛�uv]�� q��4G���It�򍝿n�9��W�Ȝ�Z̔�h{�6��kڶ"�Q����F}���xso�Q$�bJ��o7�3R	��X�@����GA�"���T��-��5�a�NOY��&�ѷv?4;5��Gag,�(3��	�M���E{Zl<zF��ň	j�1=v��Q��Ru���p~R��4Xd�V�zҒV 4C2{����X4�α�b�[}�$��-�\x���OZ�xcʥ��萒�d��9T�zN�X��|��;�0�d"-o�d�b䍙�j6:o� $e�W��уo(�]Pr�@>t�T��v���L4R�)�wdr@�_2
c��12y-�"	}��$@�'ޝ�!(��w����)QGˈ��@��[�:i=�p���IQDb����I��j���iR�Ϳ�V���!ra��N���	���� P�7�)�Q�����ac�l�-�����E�L�9��<g���by��y�i�!��zO}����p�P ���v@�'����P�$VF1us@A�ք���|�J�jG�X�^����0'�SO�Wײ>���a���	�D7>dT��2�x1ࡻ
��J6�S��'�P#�wX�`g6F�8��c,Ā.`���H��Zge<�:7b��������ᯌ�+dI~�d��]����'��,�f%ןސ�_�#��>�W��2/����Z���2��u��5g�ci��������*Q�	�*��$!t4�~M����5�J�ϓ�?E7��:��`Xhj����߄u��+���NP���S����U�S7rg¬���Ͼz���5�U�w���Vo��Y�Q���:O}=B|=y�Cm�[�y0��Ҍ��O1&����3��6k�A��h�_�����Q��bCIzN�8�E�����B��P _'���\Cg��$���⃦�����W,�3u�œ�`��u	t5��Y�*�X(�q��y]P!o�wL>��*���|��_p���@����.k.Ӡh��quf�jsQ��8`2��Q��C�O*kz�e�<oF�5lx��E_�×�����`�2�kc�3R��F���#���^hrF��֥�u��RGp�P�X�����6�Yy�|���X��-�I�U�0�v-��n�c#� ������{��IU��>��H��=<�`8B��6آ_������,�2��u0d]�	���q��KKMB	I���Qj�$U��S�:x�����C�}W����@�@� /Ir��j�7����4N0���[P:3����c3S|�4���%,_����x��
M�8NB�m\W�凉��;GLCf��N�$��Bw:r0G�Wy�{��#>����g:d�w\�hP�aC�M���[�s�^��u��>���Bâ44�4:�u/x�����ܞ�
�$75��I�:��[�[�#�Aɇ>���u ��<�9�m�+�c�bkH-��!r�r>�@�="}X�����:�C�������b}^�PTݞ��ysiͶ\W鶻A���z<�.��!q���nJeﴄgF��7��DN�9�`f�P���B%�����%���,:,=���uV89�
[�F�J�ű�z���T��ܻ���#��f���Jn�"�<4+<�Aw�i��k�/I��랣�r�V0��P�]�ylb�1N�A����>�kK���$}�Kˊx\ڪ5�_ase_��Ķ/{�#�ٲ�b�G���f�)g,�e���'ON���_�����~F ��>���@d���(f
)	�Q>L
O	���b3�'^�~I}���R����7�S�J���-Oׇ��r�PR2:�MʛxDu3�G�R�</}��ɕ֦��̲��~�|n��~WE�������ަ�Y���k��l��L�EaU2�W�k�p����+3��բ�FdU�����꣔{#��k�7*7�0�:f|� �3���F�U���� ��fM�m}�a׾o��� �g�c���{04��;y__�""ppxYe����9+=�2��%�c��8ފ����Vv�i��ͼw�Ć��z��){�@[k���K�5z��m���9R���� �i�0�V��2����7*Q��H7q.�&Uq"� �Mo�_�y�s!��^0Z�hZ�s��eԩ�,�{٣��Gt���oF9�'1cm���D���o�A�ě�g[Ca��KCrd��}R��v�f��«ܞ� �``�q����h�q;DB��wx/��;/�
��C�5�J��W��h'�Iiqu@���*�)�n2��Ge����_$U���xp6#f\��&�3	�3�ЩsY��8J��C�u���-��SKό؀b�B�߃�W�>wۺ�8ț�_f9ųTk+ܥ����y���G<��3���p>�Bb�&2v�E���	W��sy�e�B��S��sK�����(n��#��e���HiZ.�h*o��c0EU(!�g-�D6K�g(W���eQB��y-��2�U�aJIE�.'��jj[!`n<(�j&OXN~��������"V�oa�,�ы�/�%y�>��{I�r�&K��95���60�{��|a�4�)>t�0k.��Fԇ�9���s�V@���Z}������M�Q1P+Bŵ0	">����o���rg{k���p�3�p�:qk��uÙ0����c(*�ި�%۸��q�k�R�r��"-?>�sA�<h�ۚ��N'r�M���������u�j�PKFK &i�V�9ʏ4�:�r�a�]F쌆���a�]<u�6VC����-7�Y/	"�!g-�<v7�$�����u��"?<1��Pso�Ի]ĂEf:�)��H��7��M��qt
��Vv�zUMmC�cǁ��Ng��?RL�;.���"$����w�

��Jj�Z
�b�s
������ʌ�a�|5TUt��� �p��2p�iE����x�Q������/Lju��^)s����WW�3T3գ<>����u���W���"�[�i���[��(�cp3gVh��6���B'��"J�k�o��&p�Sa���?e3Okf�Tʂ#ˇ��Π�v~�up��� �YsO��"��fL*~�=E�[�|b��Ĩ����k0es��@;�1L�դ���#,mkF�*�ϻKs�	|� �F<��u�:�>	$p%�]�^�oa��?"��~>�6��h�s������MD*�9$'q2�Z��;�� \�pSɅGݭ
lB�_9�6��8�dW�#K��*��ڵ�~���N��z��P���\-6'�OC��'�K؄�Q��^o�j�]M!�<<Cѱ#%�7Ut���rA���J�PmyK��^��#j��ם�����,�9���Q��~��lҙZ9K�m��-ͯ���OdLok�%�Ì=�	�7�`!�����^VnՐ;��ĦX�������J7g��-�d��.6��5���0��g*���;o����T˒��9,ڭj�%8��B�U�f���p!�I�P ��j?cE���'t�9
p%zB,2;�P|`�L���@���zQZ_�#��a���G���Yj:���:��t��?�8@^\H��m~�zV��S����{�l����E�{���	RD��	ި��T��7�����]�����v��}�!�b���@�6�\���Z��Dc�Q��4��|0$��ܴ�̄���-��F�ݕu��Hx�@Z����op�����s�w:�F�n,�������|�x���/J�CS�ۃ9�ہ�g�,�u���wm��U�u�Cy.�Q����J��b���Cϴ�v�</�b�z�I��T\���/1��
�� ��r���c���Q�������A%}���-�7\2%~��b8���lm"��j`�- ~lY�0A��h�<��6Io�u8���lT$`���Ǎ�'���dnj/���y����*��?T$&����O���3lG)��DK>���-xo@�>�W�0��j2�YH̡M�FO�[>�B�=���6H E�=��fy��)���]DJ5����5ws�G�WY�U��\.����	~��
o����U8T��+z�a� ��Y��O��B�;����?��"��g@�i�ǚc�� � ���	s��9?�7
���NU�ʉ����>�a�iZFsY8��s��آ`C3s|{W��^�k���Ã^ߵfe�?q<���јn#o���+'A�T���f����&j�$���_FO�n\�f��ht�l�{V4>$m1���󣬃��|����G���U��m��Yk2w.�R��q{�4�m;�^a�n�UD�Լ��b���𶄦Mފ����Lw6hP5 
Mi��=T�6A��r{gl���V��e;��	�o�Bc�[�F�R�Go˼���V��R��{�0��n�)ܤ���%��_�:��Ӂ�}��L��^$c��M�\�}�d;�����ӬH�J1ƮT��ȭ�����c�k�(�-��9�U�O����%�QOJ0PGH��/��`ĤG�n�����~F�?���w�uSl�_��(-o3� ��cTi�[���'?[��d��@Q���ǘ:�O�Hͤ�{#x����������NX�z�sfaK'ǿFWH�4�[�j��Q��������&�ơ�>D�Z������B�@�0o([�<�~���p-|㲷ʺ��xzۨV|��v�4
%@��eQ5�w�$i�~�hR�uft'_~�Q�(��!N�A�q��n�G��a�R�?!�q�8��#L���=V8�6-'3a<��v�m�H���]�f�lP���!�,Q|��`���ۉ���1�k%K�
g
�g��M�@��=�󝠱(P���Y>��6r��[��.��uY՘a
�s�f���dvn����ϙ<�L!	�^�����=b��;��g�o���a�����^	g;�/N�Q�6imp������<h��ǭ�8>���o7�x9���$kdc_k���% Ca�K���m�"�ÖG.d�~NM��P�.����L�oS$�e��#�-�������"�$e�~�+�>����%I�X:�sq �K1`;�����;<�<D��r�>�Z��l$5�tz�QOZl!�w� !@k�~��	����݊H@�M�i�^��i������ ���A��J��S��cO�<�>B������S�_~��ui=�9#�)~V~2�y��>8��U��eaP���Cw��I����Z "����0{́J�u�G[���?��Y�������.K���1���JT���� �NJ�lzаNɷ�p�������^�\��*GK��?k�4�Ec����u�r���8L���b��	9�2�9�f�	��uBBs��
4I�t.���9�=*[�t�Sr��d�UVVt���� <
ޯ���O�����3� ��+袘����;Ɵ�zT?�v��[t�jRLtB[`�����(+6�F�Zo�lA�wI*i�ߔr�r���z	~3�^6i?�h������Di�s�zg;�����c�<kZ��zM�qr��aE� ��#wom�`q��n��/@�J[ظ�U��ѷa!�.[ ���!,|}��׍�j���=�DŜ!�Z`�&Qj������D!�d�{�*=�On�Q�q�T4�6��w�����V%�b�.)�1�=��FmÄ�3�N?����'�`�9����6nG�q?���4!(�q�Me�[H��u�V`W���S���S�~3*�ֱ��|a3��C�c�B}�Tً�cU���R5��Y��q%Zf4���#@#�n�v��!����D२{+u�@7�Jp�j	2�a4�%���n+x�G��:=e�|sK��1:�$Y$��?�tL
�L;{}!��e?�����t��2rl��<�Xq��|ŧ<���	��Am���r�˶QҚ��3�u���x�D�9��t,𰄸�q���.��v�7�]�'b�Z�n�Fgq���t�1�x�x�d w�H���p!v�W�Go�h��3�2�vT�}kuF`���oc`�sˌ���cCZ�%��~H�}���謑��������z/���E-�Q�瞗uS_���Us��ʋ�ƖG\
����´�X~���$�h��;��if�
�_�	�>\�v�=�҅5�n�2����0_fg�y̤W<�I?�V��r-W[��X�&w�#H�rI��_�����Y��v�e6��������'�HН�s# �d�bM0؀�p>��T�o���UR����Sy8v�SF�o������G����~�j:V^�a��m�|_(/V���f�[n�y�~4��O�%Sg��ˣK�����Z�u�H�R@�ddwII�_a7�i���֑��/�`��3t�)0�R��F���Q$g �Ƶ�/�pw>���(vd�_,��Avd}�%��7�)P��N�I�J�.o�F��MW�'�}����|���i{a�M����#�"y���*M=��@��ѣk�~��0CT��ɸ��F���'��D���pT�iV��G�j�I�;��������a.��#f��?�o�(E�&�]��1�z.�fs�����^Vë�ہ�:��+�ve	��j�h}�gѭOd�<w��"�����	d��!�nϽ��DC��{�0�f������П���M��Cd�����DXX����a3���}�7�x������[��ߧ���Y�gu�<(��Ư��LaG�g7q��=��#6*a q��3�+��ao��c����&��5�����]����8�:Q�6ˡ.�36�-�$9���,�C�Y�Q�$��?k�s7������Nm���uGђ�z#v[w�08���.b���B��8�` �K�a{�\���ǅ�>��z��rL+IO�m!a|�\T��P���_���o=i��.BC2=���x�mv�E���l#.�B8��F��i�\�@Z�����d(h�QW�B���f�@�]�)Y�-ٖf)�!�V����|������@�I��/U&X_6M��Q+��Y����}�6���R�ᯤ�}�[W�,��"�T�,�D5�ΖA��� _A�u�F�[+
x��@�:-�t����J<�trz�*��Y�D�I�^�L3�v"��M�e#\Ψn�;����K�¯Vt�2ʹQu���_�n	Q��d��>Ю�i�k�V�0�3�k^t�"��"��˻�b�p���0�i���2f!]�`$Yf��_�ѕd���
9���R}���è6"f<J����ݙ�IW��%,*�-�a�ޖn��+.�����뼪ڽ��缬|�3�}��骀����&v��߳x;S�e�R��]0f ������Q 5@��ƙ�f!1ђ�٠B�?nu#Q̈́�*Ӗ���
�u�m8A�EL_
�>���
"�UЙ��V���Ʋ���].�"iy�*jknsdw�7=�㖕�����foC�@h+=�r�GCG{:�4fZ�.�p�7�!�y��s��u�m*�E���9��7?�7��}~��Y����O>�_(P˧*p~q���=��&­|`����D~�ڀ������R�-�N�KNt��(�̦;RG�Ԏ�N��P@��"ۦ�>������k��֮��(:��v��Q��&�R��=Wl̇�f���"r�~�n��.�z��!�������H��e�3�΃�BZtP,`��W�sICjNT��fzq01ѫ���W�^��"���~�nQ:F?��j8
�5��g-������?H1G8P�$�Ct=O�uv��ۢ�mK��ގ_S���j��'yӣ]���D�,S�gNM/B _#�ݷ����Շ�SI*J��$Ap�wˋ����%w��i�kbm��� _���Ip�φ���j�c~qs����E�����O��{e��t7�] �D]����p��a@�b��!(ڤN_�٣$q���^T\~��'q�	�l���9}���P5[/^��D��	���T�3��1JsEm{���dCW�W��;����E���g���De���W�^�8Oƹ�}�O�|�/��dc�2:���o��m_C�*�;����aV�u�|Q1P�[��)��6�'B=�����bi�#LzZ���Q��K�I	�mWj����Jí<_m�{_Tg+OӦ\�z���䌒���xr�MXG�5��$��)�pE�0�ީ�o��O��2a�� �,�A�\9��}=�)t�K)'�k��[�V{7bU1q�nT�C�C�k�廣��0��0��`��� �	�ǀ$y{��M' BWi��T�n^�j���i�8�!��ݥ�H�J�tj~����/��B�I�f���4czwl��`��ډ]������*��'���xbJ�*��j��t�CE���N��6�/9�����y�N���^��x�y�V������'��E��������m����r�<�Ė�G�m�[���������9�}�����ի��Q+I�o" �u{՚%��/K�C�_Uٞ_�kVl�c[kC�`M����?���r\럲�d[� �=�����ц�<׌*"Ѽ���b[�!8�}��4�i�
f��?�Γ��Y��~M� ��|�W��t��8t�H�����!���"�4]g�b�y�l�z�U�X#uSO�%�z�٤���i"�_�(zHé �Cx�����a����Bxz�V�״��LVА�����4oa&�t�d�q���`,X�u=�����1�Ml8T�^6�>�K������Kp��:v[ֈ{�����OEj�e��<H���ۉ*�f���GPNQ0��L����J GV��Ö����b7p|�s\��u�C�vS�p��kL�"��.�ň$j�V�[r0Q����hR��vU<�b����qU� \L:d���a�z��[�A�$A�
�v�a����+)ծ���iy��9�@f|��%yDW:q�5����^���!���]w��\���� �×���a8a"�ą3c���[}ٯ�e�_9�D�^�j\˱�E �!cS�A�i?��N���0��!S�JϸC��@�K��$�B��+|Vȩ�ڢ�0Y�8�n	DP9�o����������,{l/$It�&H�o�R�D�1t�S�>I-2�����	��Y�鈱��(��炌�ĤlB�o�],փS/��|��:��VT���1��� W�<�����Μu��/�6��gk�aj�y^RY��шȦ e������H��#o��"���AH%�C��<HQm�&G=�P,�l�Yw���H<	{[�GАA╿���f��r�/�~��Ƚ� _��j�1N!��a��'�㰮ӌ[�;�y����&.;�'����-+����6���|��5��^$�ؔǫtJz@�*|���_��O�A ������)*<��\>;u+��qe�1��m�u�d�k;�����uo�EƳ�sK�$s杶n�P�2����%�]s����ؔ�����!l��u��<����aY3����O]��V�Ӫ�P�T�M:�>����v6��)W�`#Fu�0v�2�2���y\�����x�蓮 ��U2c�{µ@�8�l���S���0E�l�6�_��E��/�UR��lJ��ɢ1�P ]�5mF�_čw��߹�~�����`��4�7+J�:-
]���3�����!W��ÝR���Z<ༀ�Z0�D����_*Ma���1�ie�����T_���������h�g��3�7�I����[�W>�����!�<���vU���P�'ࣩ�Q������]���l�)	�>��M����8�%/�D���f� �`�3D�>P�R�.|Fc��zO�훁��ΥEE2y�����ɷ2����PPP�s[��V�eQF�r���V9��{H7���y��
�vP����9�O�:}}	����J�KW?K9��~��2{LL~'�^�S��C �J�r�Ɖ�,� T?�!t���I�|�%����m.\k/eŒ#~F���j&.ƀ7����Pf�fF��>uc ^���1>��t0L�Қ��l��O+2�M��|{8�D5���Vse�۴HS�P����G/L��_��\�}��-+�Mn�s�{�e�!�9����Y|i�K��״ �+�&��z�H�>}�,�i��޺.�b {��a��Q	��pն٫���9Z�i*K�Z[���� �'�=�癩gҜ�u��a.�}�hv9Unwܳ�������tqt���ډ��V���6��|���F�Uû��ݗP]��ԙ��Rp-������o��g�����;m 24�������ٯkD�S�|w����>��A	&�����Z���Z��  �2w$:Y���\!oH���5�΃A�[�s`�C��q�w{۬� HvIi_#k�.;�Q��3U�8�xD�)_/��Y�W��'��%�/rJ]�Wr^10�f����\Zs����=�GT��e��%�ۀ!�qX} ���k ����&��'�1�r�?M����S�%�$����@f�	�$���Ω���#�],����X;�P����Ň�$��V�����n��