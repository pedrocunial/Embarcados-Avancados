��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cЌE���MuW�H��I��~�qf7B�y�g?�:	nYg��-��~	�c��j���@3ۀ���=�1���K2/�e����ׇ���_��틮! O�}رH�$�n�G_/�o�d�+�`�������&�S3�q�&�{��B�Ӻ�>cY�Q=�"H�q#uDܯ>����7x�w)�xӴ�u��O��dâ�sG��R��"PY�
�w��D�[��T���s]���_�(6��b�x�j3��I�����V�N�m���>�,���5 �#�ĝ����B)��:[�\g���nxLH�wS�5U\?(�[{��M^vﱔm=���$	(�`�F8�ZB��A@�xkj��|�5HA�]�D�V#�|�����I���S��3$�H�n�!4�p�V��`�4mXT�?����h#Y���v�P^�* <���l0��}�Q]���M�t���(�\��N�ʳL7����Y��U�Y�!�!=T
َ�T���X�k�C�s|f]V�<=�%�s��G_�I�m� ݤ�>ܦ����pL��K~z���yf�N��g��+$���秆3eT�=���~2�e� �u^<���}�4���AdEsv=�磊��ٺe��7vN���q��x��o�W���������Q�k9 �CLT��ei^�SsO6	����}�S�ʋ^xT��<�P�}�-��_؁�"��T��U
�@f1>Pn_ �3"����A9e���T|����E��I�o�#\39+��Fl����LE����#��r?Sl�kk�o'<�{f���d�0�B~it�&nrj�}@��x ��_q�&ZC�����ӿ``�0i��/5���[���V�e�+�,��1I���Z��ׁ�v���mqLO��4�,l��=y�f���"J�0�TN���3�bM��]����v����'�ڎ^?<��#�S��3��-��osH�0)B�帚E,�䕼�<7[(�LXO^C/[�H�)үd�|�=ạ��*>]��ŝ�� ;>�ldyO�"�Y��� �H�Y�*Ҹ�R�)3C�<� �xu�r_�u'��9W���T���AƔ�����r��B*΁�1<Wn��� �OM���l�0��¦M�I[f)�i	�w�E܄�O%��nbg�d�c|��Ym��o�1x��0�x�������q��cy�f����J����K�8Gdޏ
_f�! S�foi4�Q�������Mj�	��&vu�V �~���^��l� �Y�<ay�8%������)��tV:Y�i�'��~m�8��GVU �� G���OTu9����)uVzP!Z��O����B�{�(9�l��� ��t�=��
��E��!J�}���6}��x룛Ҫ��1-Q�hID��N��֡*����p�5��=m�B�zP�?U�uID�
�L�U���u���c��?���{i����cD��c����Ĵc����T�w\Wq�?6K��W��yMh[�`I��kVB�D�Zܗ�xZ������H��,��X-Q��Ա|���6����t��Tr{-5[��c*^��ݥA�`3u��י��0q��{���6?=*���-�U&ct�@9��Sn
�5�X��п���")R��֘�U�R��,���6���w�UI�����5n�s�4��y/�*[���S� (q �q�g��Cܼ���u��#�L���;�4���o�݋�y��Jӄ��s�3���p��_y���k�q��f��ˏ�@5��13^��i���r�6��C�Go��Ӑ��מ�7˼w��a��}8�!Gzs��2PQ7��;*<~ ��".s{��\7��H�t%5N$�o�A��yS��}��`�"0��g��v��.�&�웼8㘈No�J��?j�b:/ϥ�=Lk�i	Ǌ.�����G��_�r�n }�l��X�ͦ���y�^t�T�ɬ��O���_T�1X#�tX��0��3�F,<;��]�!J��U��g�̮���=�z_�+C�0�1i`�:�n��.���9&�0�'5Z�A�z8R� �7d:t���Q��)B��5UG>��
�i������`<& U�!i�,�z����Y��ep�!6�A<�\R�	˨�3,+U͵*b��e���>��k��^�Q��{����T܂��v����T%bJ�U�>��P�ۿ� ��!BgDH{�k���*�'=X*4����s���8�OJ̩&H��8�=��Γ't�=�u�Ӭ�1�c���Չd��[S&�\�Gd6@�hL]�	8�^�V�|��J8�q<Jn�צ~�>�T�t֫��J��=F�]��|4�f�_^i��C��C��/��c�Ϲ��J\ts�l�.��A�+��������[�= ��u�l�lJ��Tc���0{ nR&�*B
dF��Lqg6�s�.�WW�����
I��巙�o �������b������ ;�b��Y�}�^&4:/!�*^���F�Ψ�*f�p�'�i�R�ۜ�.Amݐ4鏶`�^�2���spy�����[�����*v�s7$7�(�9�pb��۱Z��䊶�w�i�Co�7���x4����dg�5Ҿ"��I�2!8>T�D�^TM�#�d�m�C���_�$0z5N��͈�b����7V#���6���+��'�֥�o����?T�QUe�`67[�A3������<j�����]4R���;�-V໱��~���<�1u%F�2�y\l�jZ:iΏDcQY'��e�9�#4[M���"��"z?r��t���P�x����M����pcr�J����5� 1��>,n��������x {�̛0�;4�	��z@�m�T��wCc���u���X �;Co\B�5u�PW|��k��Il�!�K<w�RH�?w�J��4�3B}X񾍿R"hpQ�"^�5��NM70d���2��D
�}��H��$
I��{Ca��å�=Rʔ�`��QV�@���':c��q�u�3��VZ�0�!D�(	�;����r�	��YD����\��\	� �!�C'��+, Od����t�2s�C�}��� �"��Xw��&A϶TϽ�|,lb�{���v0gª��%KŰ{�J�^�72�V1�{K������r�OZ4�ɛS�_�1�?@k)�ӝ�~uN�b��E�;)h�Y+d%��Jع����|u�v=�z �`��B��^Pb�>�ٯ��1a�P?��U �ExJ6pQ�іx�����e��譲��2[*<f���dc����]=7������­�o�m~j��(��)��OMUG�?M1$�H��'8_/�gtR�~r�|7�䍪s_��Hx�>0�a+m�5jN��<1���������C�~1�p��!�w���z�e���/�уCXϦx+;�*t���cp�)gN�%^uu/��?����j�@�1�Np��!;Ҝ�2���~-��߁�9Y��e��$�&�bk|ܓ~���i���X��0S��� ��9��n!��f�bz�ʄ!sG,u��P�z7Vm��(sැZ�,�/J5K��޶�w��@�M��A��~�=�Ǎ�����^�d;��(���F��0���#�1X��o"���j��>�T'��S젝(���/#ǲ���?�č��3�؋�<_� 3-�lQ��:qث�8ӯ���@�l�g�$�NGNϿ���j��7_���5^���@��w��U�_K�l�A��G�{e���
!NWJr�+�C��������j6Y�+q��oܝ� (�Lwahh %]����>z0�Q�\c9Oy�S�i/+�[������ ��<��_#J�őn,�,)�l��Ď����k�a����� d�l&g��5Nw������dR:]b��K���U	XH�� �*�dK���[�X��;`���G���~���:X��A#̧yU��}c�} zN�J@��,�՞4�s���Kfu�M�u�W�\�[l����:�1!^#�=�ұ"ץ�"��KB!:ƍ5t�mq��-��$�:�؇���EM6�͘�Mm�,���ɨ�Xp�����bW�u4ƝvB#��E��~~��HT �Q����à�n�� *��&���־��Ҥq ������.ˏ�
3�X�P-!�b�I2T��%�RMfi@�XA�v��\'*��p	d� !eTd_q�` Y���q��s�AM{.@k�}�����X��:>�ݞh�����EG�Y9}����"nvDPzF!VC"|�n�W��:��d�צ�.8?���x."����mZ����gCE�G�Sxx{i���e6|ܷ%>���4%,q��06��V͟zc����o��l��Ӏ�����Sz�n'-�^{�i�hQ���u����凤�AꆾС�K�y]�~�N�s�T~A�Vx��7��w�rT^�`��h<N	�bց� �E^�
��x}��4�	a�n/����G0v� a������IJ�;�x�|��d�܊Y�W��&x
�C�+x�l�)�SOWI������M�[�ֲw=}�t\�HiZ���XNBM�@�C���qSQ��Ot�P��L��r��e"Rivi���d�j�$ն~]� l�ڋ�a(_XFf���%�3X�QP���\8�.�sw���R����{���r��O� �AU����a�����c�۷'xR�Ē.Zk>����^��T3/��> �^^�ow4~�_�c$q�����p�(�uʶ�<��6�o���}� ;g�z*�i]m�����	�0F"��2/Qi���J�Gׯ%b�T�c�}�D�ɔ�#p<HŽ�?��
�G.p��Fl\�L=������		�('*t��+E9+�e�� \ �;K������hZ�>�%$�F�liM����a6�0���8�`}?��r�{��_9�z�A"Ew~��%���{EC�#���C{� ���?ƣa��E�g���V��& �eb��{��e# �|�`�3x�.ؗӥ�Bld����'�]f���M����}��!ͦ�$���Fh��5��ꠥ��U���KKR�
p�&�N*�[���Gz	U�(���F��^�<��k5�$�L���8����<b[J�9C�{	�����4�:{���X��`-\��r����t�I����������@}�$30i0�8��F�֜��r�FRZKBp��͏2�߲ʞ�`�WH�D���ׁ?7�xq�k��dh�S����,W��/l��g��c����s�їTT�9�Z�s�>�O�����-?�ÍL��Hz9e.��vrь%�o�Mx�E�\���ܴ(���y� ��MY��hݑme�s�`0z	��#�e�.�S���R��u� ��j������2�<�h�2�+IydV�u6Ag!�I(�k�owm
������]︞�U9�-M.��	T�u�4o�:\9�mF[��"�<��,�|� ����N����ۻ�g腶k�wڵ�"WIGJU���������[�'H�'�C�	~��_/�~'�^w�~�'�4u�aY�v�������j���*>Y�;� ���3�ȸ��}|�SK��L@?����i����t0XA)��pW`~�� ;��4��G��?
����oرuv�c��/k'q�$`���0����ПtHUg*&��+��l��b�z��ӟ[��1��H�1)�^���fMv�9,|��l���oq�R�ĥ��:a�"
����r�����ő���p����,!M�ˤ�����B�_L��WbZ���2�샫�Ɇz����w:�Oq����C�������Q6�7��Mvȃ�rТ��AQ��Z��Cr�!5" x��-�k�g@�c�G�_u�j�_&RLS�����W���=$J

���/���W�=�1}L������:����)��z��#��E��_*��j�?k���У��jF
�c�Z���U�R�i�<b*�$�e��ZZָ~�����3.��6��:�z���#]@�^pԌ���
1��B�?�Еs`̉�['B�,�+h'����J\�Hnlx1���H�8�=>��/.]'`��R��3ze��%I����
g3 ҏD�t��@Ʋ��v_.L�?�w.DQ'���7��4:�$zo
�z�	-�H��L�\���-��àQ|}��J(�Y��KI'qG(~9Nv��WWyl^m� ��{=K���x~@�l��c.�I�Qjz���`����w��iƤSރOd��]����l��܆�����ˍ���e���x�]�c!�E}�^��y�7��aF���x�1��I����g��C �`*�V��N~J��o4�E��s_��z��A�ت6��нrl <�a�@4���jn�w���d���Q�w]�wO1�~h�7#O	�#A�
��6���@�Agl^��^����Yp�x��`l*��]Z4�.���2�AR�C2(-��8&�1�����8�T%��j���v;y$�������Ą� S�t��Co�X�D��s8���JM��J$���Sqv��siΖ�"fk�[۰�5С-D9�`�������$/5{� H��}-�hp.�p�C�AT�PY�|��m�Y�M����z��I�^x5�@���-?���
�Elc���K0�Ғ�Q��C&��A���F�%������K`, nJ��Fj	.��~9�����7/{A���D~	�^�����#��k������Wt\��|����2b�R��3Y�X��� �xhW�O,l��3��j� �@%'{#���!��]��� ���U��N(n.v�=z���qW���@׶Jى.X)���e�=��bUA��E����CQ�~&c�
E�!�(l�F���B��h�Ch���W4W� r��3���{\�x�V��rK�A�����=D�D��F�����4���v�.^@ �9���2[�wI��#>�oV/�+���gzb�=+E>���ޤ��c޶'�D�=!xo�Pg3]s�A�B��0���C�?�Q��1A�L���bU���A"�S]�ǻ,�2A��_R�5.O�I��S����i��L�2�;�M&��喛�D�}�#&��FV�+j�q�?w������?U�
~�9A&rXٚ��٠%)7�[�p;a2mV<��x{�T��W�-�"�GV��D<�dm��g�d���~}��ؼSt�^	ծ��f�����
��OU� ;�qb�/�)�����Ct#�S��0\��`��mYb�6�ɷ�{�\lOm��������f%���
^*�)�j���\h�Ń�j�rܗpL�������J�1x~qܼ%��u���>��u��S����f���/���������T1��u1(H��N��$V_�
�g5��*�>�δ�~�6�oך��'��V;�����ݤ���_�uQ�����<Z������������=�#���V9	w����Y�7��������L���޿(!��3<���6�c�%gE|����Y�$�'Ô⧀
f>vk.�O@Q�Y��N#��&��Z����ӽr��d���Ojѣ����P�'���7IL�D[ip���c���:�Y�q�R:��b��Q��ʌux6�\K\�P�;Y10^�_�|�,�ku�碑� ��2:L�U�wşg�=J�\4
�g�^~*C˸����%�y��QX$�R�+�=�epxYIU��t����_����~,F�J	>�K�~��� ����,��ꄪn�	�j`
İ��#z�q=�?��g�>6���BD��x��ǥ�`��H�2�f����9A@.���3*���ZGXf�yj��!qd���d����֮��u��V�%mK�Z��T��2������;�f��:�\��*���͕��=�H�Sv��@e�B�L��;&��+nJ�!_������g=_@����as]s��qٲiYVv4�@��6�н��ǣ̼�_q��Y�7/��N΃_��_܅���=���P��|��@�g����	*;����\:ڵ\b��VU���x�"�l~�+�m������sQ�����s��[���H'�Z�����V�_�k��~�Z����ltc��%#?�m���꯯'��S���䬖o{*�f�e@ʞ�Q�n	P6H��b��@hϡ��=��4��b���>�2v0:��"^��l1�'A���~)�|FZ;fUU���Ot�17ڼe�'��<ND��(�M���ֆ��o��t��C��~
~�6�k�V��n���~~.���/� �����K(k?�D�Q��t�.�� �M�����F��.�cw�6��pK��LV� ���������,����b���=T1t�������}7�������\kGt	w.�Jޤ��'�<�։̛-�:q0����]Gm�ΙW�7'���:������|ka�5���*�߉�A]W�"<!(��m)���{a��&X(f}> ��B�&�p��j����rԟ��	F˜���΂��$�g����)��PzU��~�'��6�X� �e6 �487'�F}�r��� ]k����N�qLb��E+|5�Ȳh�����'S�pඳ9\C;>�#��F��Ђ��M�A�������U��wB����Yڝ�H~�z��݈�����>v�g�.��=�~�I	��*�{���i�MZ�݁0x?�z�翑�Sq���	�{����o�;�7�21G2��`�aH�L��}�2�W�FY�Z�4Ҕ/z��J����_[�S�.6Q��,X ^��Z��z^|Cgw!q�U�Z���KK���cb�d����Rs�˄^/�v��7���\|	��[��\4�J�W:���v�eok!��<�4v
'D2�V�̟�B�-3bC�vY���PzI�cb�v�`$�>vˮ�ӘI�	
���,I;�n��,y�w K��
b|�S���)�(l�<��~GAAv���m�*X�ѫ:��������p���H��KEp�������T�SUa������߳�>�@��>���0z��[Y5��t�n?W�;�jG�s�lBǴB���zG�� e �y��F��}��žP!���y���c+1�*���hB��kG}�p���z|��ф���~�b�e��}ǬD���f��"���q�=M�$���� ��##,xD[��� ����b�µN��ٻ���E��?{�E9��n;Ͻ%�3��.�0��P��$$�Z��]���"�6q���S�4&5#��/+���Q�ϯ�SN�{� '�G�"6��L۞M�H��)�����MyP�=���xL��&x�#��l}�H����1Z�z�m���R܁Am�}w;?���E��ӮB޻mei{�M���S�d����迀Yf��mՊ�_�8�W-S�R�o.�4�+��ӗ;�,���<J�	��mEow,�9���\v(H�n^J�� �s*�^� :R�8��x�,�If�Y.YD}��Wk�*�T�(��d�i�j�<�^��w�C��.Q{�߷�)����U)Ğg<���H-s���N�EsQ<�m$|�ºUp��p�s�Ԙ\,�/��PB���2P�J�D$�һIiZ�o13{�㒭x�t�_�&�>�sn�d]���2{���̼f��li����)���_�2$���	o�e��iE����5_��/�?�T}��01�2I5�f�:��x���A]�g���f�ު�}��85����a]u���\#��M�� �i��lI<��PZ���0We�2��<5 ��Y�-�;����z����fuju���I������\e*�:�V�g�
�>V?=*A�\�*?8k6Ё�ۗH
� �mI�Uŗ�/�)i���"�Ft�j+c�#���C'��T�5_w ?�R�N^ ��j�͹H3U��9�Ӕ�����?����śj�Xt[��%�c��Q��s�´�uX�:�?�H��Fp?]�uzi\7�\!�!�5��G']�Wd����|6n��Rl�zoŜ�N��w��6� �����v@�{�}x�a8�"�c@[UX���OcC�x��ѭ�{]OJ+y�;e��\5ؐD��б�}:#$�G?��=��/�2'��zCN�����R�������ՙ�_�^���e�(uS���Z�"�:�^ފ�R(�؄ll�"{}:���y���[��i]	/2�7�Guh�]`�;8�7�E]2�t�/4�e�c��}���c��b	�,[ �?6�JPfݨGc��#��0��@(����%�?_Y�T�=rk�jf�>L��.!�R�X��i�3|�m�����w��18��Ó��>+%d(y���k7h�J�g-Wҩ��p�u�d(�T��,q`0���,�U�v���� F�e���!�!���nl�J�Y�ϋ<��	�[��d�&��L��sy)��L{����v�e��!��Yl�N�³{9y�v���@���ǯ�猰�����˧����uУ�	�+�n�`�%�-i��m
A
�C��Pk�c6̻� V��m`Q�}z`���<������
��U6�����ޙx#1s�� �`-P�1
�Ssp�{ú�i�b�0�Ӹ�� R{�诐�i���
j��~�k"�7�O�$���_�ҧ�~IPHʄ�Xb5�$2�U���+ �V>U�!�:�k��8���������k�j(e���ʕ�������?xs��@w���Y' �ܜa,ʄ�Ȗlx����<���j���t~4[ߵe���Bm�}��yԥ���!y�dDI�W���,�����@ȱk��JQ�@��ȡ����+8�/Q ����3i�p������:h��T{_�n"�",�5��۴َ�Q`��Ŀ�J�E��6�G�'ΖW	Av����M�t�Hv�ƽՒj6�}`��,hl&�hԴ�y��'�k���퐿�\>�l���£�JS�r�%��]�T&0�.PZPW�)H��j}�'�d!Z�g�I��/���X|�ް��E�d�8�m�|>�����{�}cqEI��IlM��($���O�Q������ȱ�=��Tlv;����N:�5�'�ݗt�]���EN`�W3���;��1�,��N�n�J5�Y_��/9��)r��:bl/�S��v|eY�����y*֎;��^�@p-(��:��X�nʴ����o!z|��ļ~����%�>��G4���.ݢJ��a�����~cVU���6��.�)a����ȕl���!Y�gT��m�-��}�D���6���f�2L}�8��g��wk��,N?���7ۥ�]ϰ�֊E�ST���Ig�� ˼�� ~p	�+*��ng®�x�C�Y��80�V�6G (F
MI\�zO�4@SI��]�^�ǩ�O�	뙒-�R
�����Ι��8�!	��X 9��k�N��$�f[Y]�g@�e��f�c��%2�i���
#mrN�ifWo��M�W�D2Rѵm_��rB���L�[7�F�B�B�k ma��g������������HY�C�)d�2��.�V�f�������̳���j��b�v�	���&�k���n�c�R�θ:�.�a-�� z^��?u9W�YC�� �=p�4r�@��"?L�CH�kH�� )����[�f��҉����UM�($a6�H��-XfM"r�cp��.q1��鸳\�:V=���:���c,X����]j:h�+���6Y&��={���m�A�)���F�K�խ�ƆT�5����5�΅�h�9���#�;&2|N���X8q��\-�>Rii����r�$�3gaw�%��Y��1RO%�c?\���#�\���H-D�n%�o��3#)�*E�)t�o9�3M���o��{G���DJ!��F��?���J����(�v'}����>E�U�K#���|���x�&�-��ӕ4�_i���X�3���tX�.��nx�ӌ��Q�N���c�}+O�7ǹXY�"G��0Hc=��6�x� R!�����`	�:�
gt�����"�U�zS�{��.���@[�����+�o� 8�j_z�~u'`]RZ�8?K�#k��K{�����)�ʾf�i|B�����haB�S@�ǂ�)�=�%|��C��7ru,K��Q����e)MZ��������fo��)	��Z�R=���\J:�7�����t�r�4�Tʂ�t��|ľ~Z�Uz٬Dh]:���8;<r<�/�OK���G�S[��uH{5�O6���鲢��跌��+���mRҙߒ�Aj[�ڑ��Y/��}���p>ew�S�R�Ubj�'zg�~��O!��]��D��"�R^�~��(��H��GQ�˫� �2���U""�Xc�tz��Yt��ѷ@���v�Y�Ⱥ|v��ܱ$��Z Bi.�/1:q+8&[�L�7���*��M�3����酏4 �����d�4"��ֻߩh.�U���a%��yꫀ:����lNU���C�B/Qu��H�7�/��mnh�����Ɩ�~3��KhN8�a~v�y�ޏ�ER�Cj��/�z�.�]������3tZ�8٪ǻ��=ݖ��~�v���"�AR���/���x8��QC !��rtO��>	��B���{jg9?�7���_Ex0�����mѽ �XS��7���iC��H,��"�>s̋�ƾ偘�ɭ��W[a�y�7�lsl�2\\� ���頊V�����X��EA*�m��>~s'�Z;g�\�,0V�WJEzϛ��S�G�޹�����j�������_��&e%&��Q���{K+6�����-�f�h�>��]̡��%Z҅�`�7�j�C��L�y����W�ى�KW'!��/�]���Vn�ea=��P��ly+~c����6�D;S{`]����@��p�F�8�{%��%�4Sb�j��ǳx��k�U�[���Ɋ�uq�4����QL'<�C����yBu2=�Y#�Q̍�F���C���&9���	���X�F�¥.="�1[6g����N�Xm��;����ɷ%��ϯT�&F�Rv���J��� ��
���.��ť ��Y7C��b��᏿�����hAa_�js҇+W:��ȉ���l����}]��0���&�B_��t�������fTWXm��7u��)3C�����p��\��t��@N��+ک��:�T��qǏQsa�<�!nX���k(��N?�i�.V�zm���+�Ac�a��PP�BK���>DhP��?6,ӯ
�#,����yӸߝ����v�ɡ��2������2�P�u������&� �"���+�D��mD���(�:U�1��o��d����7 �H!L����QX,V�nt~�⺂��v��R;[��$j���B0qaֱ�;�Wh̄�uF���#%T���hz��D�o��=���J��0��:-��W�ý������j������Q�1�!���Fw�n��ӱ"�q���
��01^�Ix��f�|�	{#�����k�ie~q$J���Kz�!�#Ξ9�~bWUg���y�2V�h� E���i�����ls�2���T���H�q`��W��w�N;c�����	T�Fz�d�s�8��Pk���Hv�\��-E'pMQH�6�W���1�M�� ��w��y@���3�£ r8�k�Y q���}Xa��h ��C��;�SRw��wh>�+�6��)��0����Ф��i��#�\���,(uțt��K+_VL��"��ذ�k���1�h��F��h:�(�ɷc ���������
�&F`oV��K�d2o�m�!���r8_(�m�٭N�;J�@���6ODDS�w��qo'�K�j������Љ1ok�$˫���M"a���T]��\F7��