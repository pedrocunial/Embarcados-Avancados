��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c���ѢǓ2�Su���;��e� ��F!7���}�9�t�.G
���%�=;�4��#����lki��\�JG\�{2"#�	�'^����h����}(��T��bI��{s��M6�$�@߷�D��C�CAB���רQ��%�YC߅��;�<l��q��J@$n~P�3YU�=�K�r4/�lDo��'��?w6ů����w�v�O��1�s�c��7�BR�]Xo!3v5��_x˳L��3ob+��Q޹%tVl^�8�9`˵#_N,8P:�~���6�z�0��x�w��v~Y���Z���x?|>�\ָd؋��cj�W���!����lXجZ�M��������f\��Fn�_%��Ç�Dؑ��=ă"�.�ܖ'tqT�;�k�=�A
	x�G�G}m���ޖ0�]\>�7�̏(����G~p�W9t�*N�e����y(�Ȕ�C�i�����	3}�7L�i����B��Q��G_%y�Dm�S�0,�;�;�s)ˡ��=��ct�|2M��&��C�13�mͷ2'��/��ʄ��0�5�a^�2l[��p���͒�3x����>�:D�,���?����d��a�K�m�j']�����O��wB�u\2�1�O���#��F���p��?V��}z�wVf9�ߡ��w�44�|�*�GB���{җS��L�Y�LL����/��yo/���|��Յ_������%-�p��{�C��z�.͛Ӱ��V[@�0�-�`>ήփ��߂+T6"(��6�u��w�q/���`��� �����&�<z�	�D�${���SFn�RI�j쭞���?Va6@�{巜N9mk��@[ ���%)�b�n�n�*y�Q��L�Lw&�/d��V<-hm��
��n��p<܉/���u����%�����z���!Ђ�;m[��Tq�g{u:P=��d�u���(�S��4������o��c���<��O�Nf#F�ԗ�W��6�{��%�R��*���*h��׭/f�L���v���eD8��;I��6�+E���Y(��2t��_+ ��r-�4�\Q�1�|�H���)E�^�MN�UA$�e���^v1<c��	x~��yz��]Ӎ*a7n��C.I \UK
Ҁ �@�A�	P`�o�b��no�?7�Q��['~�lr��:*�x\�>L�m�}7<EZ�S�|�����#��r������t�_��V�b��٠M��h�'�A '��x(ȡ���_�#��i�QĻ�h��6��T�ٜp�Fc=�7(^Ø��ȡu�~��~vJ �T���N��������K�3�4�c�t9�+��<���ۖ�+-��.>}jj\�dE��k���A%ё��W��^],D�l����GX/�=[=,{n�}e��:�.�F�\�����������Zg4��\�㯭�I�($���įR��=ID<p��� נK.�ym��=%������T��v$-|O~,�<^�lE)D%4*������
�\v	��0���׆��$p8�|0��7����3ޒ��4\_���6�<�'}[��i�Y�y��Tӎv*67J�,�@�帡(�/�bf'��^m���X�����Wn�^�E���O���$���C1�� ��܆̖D�:CX��Чb��9�h1��R�]���
/B���K�;���h�2��f8ZQj������=�iz�=����>S �*ԉ�@�3O����7�Iz!v(����,��������a"��M��+9��4F��^P0؄sĊC^R�N����߈zQ�G	~o�o(�:	^�}}���<�6�o3W�Ԁ�so���yڨ���J�|���J��~�"�φ �go�6������%���F9�pE�[���F$4�������n�p�㢗�x�ݐ�݈�����ɯSҪR`,{�O����X�7�*��ѵ���K%�����,D��t'���DJz�ܦW���p�pmjr	+l�������+l�z�4#s�0�}P�ю/�"IwUnE�췧�y7E�xaF��g�b���nD"�ZT�iMG9"��=������Jấd�"G"K!��}W���o�\�0A{����Ϙ���/�XS�e�n`�7MK2b<�R6)E�k�����-R�clm��@��@~�F-4��ַ ����pV x���}
�1�vl)px*v�w'?�Gٛ����Y3����ɤT��_��K�1��xI�FO�+�U�ߑ�g�?.T�
f]��N�n�@�b!���WA�7�"ߞ��7�?Z��C���G�,^�!�,t�>l��'�G����f�B��[ٶT?�E#�Q��\�@Bmq/p�K	$�+F:���ʓ$1+z�uߜ��-+��W,��أR։�������]SD�r�&*-���K�z60�s�S�d�y��6S��=��#709����t����`r�m�*U��|p\tYǀ1g�^w���&��8k��pi4%�^oF�3&��ö�~�i�(���q�u�V �T����n�4�/��5ߍH��JP�r��v�3�����,6�D���*�Ҟ����4�q1��	� �9?I�x���dF\��+?��x��l� ��H��1�!&�!KlO��(3�o�s>J.QTV�*Nt�m���~���o�� �lX�v����鲊4 ]�L�L��~�tq�9Z��; �uᰫ�wL��ae��"<���Hj��0�	hm"���60h�������Ⱦ+�]��^s�@_߲�����Yq�|ǞN�k����Nzw���&���p#�����̙:�u$�2�h}����.읆.@�P��O�V����Y��m�ea俄�� ���l�>:�A�.��Fƙ�T��͌
 �v��Xl�%�8��.�A�,�1A�9|���:gΪ��x��_�.��}�����|�t��$=o̤���\���A�������-�p�|��mÓ��kg	�|U����If��aG[���IeSf�y�^Di˒FA��q��$y{�8���-�ԭ�����OH�(Ei.��L���P)Zs��ؗ��<Y���dd.s�F�&����!C��cHi�}���ds���1 ѧ����T��!>�x�H*�Y'&��YW��e����u����h{Hh�2�C*%�����ä�I�%B3��L0�|���9�(Y`�2<	��P�7�b��٨�d%;P�����á�nFN��s��d�+Ԡ.����v����H�·���(�I��4�s͝��z``�R���M��p�MînID��ڄ�N1,9�l�*v5�lΞ��ϣʔ����)_�$��
��*��O��J�J�%���@�b␥�0]�%6��p''��5GcU�}��:/ =wSx�7&���t%jvx��,��������V���er��U�Z���Uf��+{e�1�e$��8��:sw���\���W�X��� �3a���r�)�~e�a�:���{[��^I4�ݮb�>]��&�\^mV��a��9�'iRjF�z��	cI1]b�@%�Ϲ����=_R�x%� H���?Lr;��1�Dbd�sᅗ/e����&cb�h�۵�Q�Z���G�D�}e�k�o��
9�!�ap���Ak�兗��([#�͡m_Mn�y�'Y��L=�ǥ ���lqX)GQa�D �XR'BG3��!�b6;)�M�J&AiG�3ў���i���R�Q����7�:w�&̧��D�Jykp�Ԁ�S� �g �]H�ec�i��B2�c��Rf��v������:Ԋ��pj0s��#"��2�쾭��	o�h J�Ix_;;�U��.�+2�P��$gG�M���ݥ_��_��&�͖�h%}����:--�G7�r����{i���ň�)�(�|gA&iJ*�K���S�JNw3��>t��~�E��A��~%��n��V��ѫ��p��@�S&�.�cj`�M/z�����o[��jE):M���{�m����b��ܴcN�Ȫ��%���L1@��P��uF=����g![jʃ5�zF�v����\,��
9���nT6GI&�@�4A����6��!`�O�����.]
�ʧ�S.7�׉�mư2֭�M·�`Ь&��^��Rit6c�-ߩ�%[�vT����O�A �%t��^�=�V����k�%Qz��M����tnoFtG��TTt{?����8��(�/�L�Jeb2�b���bV�Tr��g�lm�s)�{�G����h!���xZw���R���s��c*>�؃_��	����m*�B��,e�K���[�;Q�Uy�$�e�#0�U�Q�� ���e�{x�~�!̧�L���4�ʧ!'-[H�V3�zY��n��93|Rzy����.�MȻ��&�f�\�S��_������|�qV��'��x��Dc�1a��H��>L�(���a����@D����q��5(�,{��,�٘9���a$S>��[&A���5����_��������4���G��&�Jh3�M�?B�}A��<���o%��e{� ��]_�*	�몠-8�1ȁ/0����	��tdf��]���xf\�c�U(�^ b��DZ�F�+}r)�sTReޡ�uQ��[�c;6"h4y)pL��dڟ|G���K������O�k���h�{��Q����a=
!	;��s����@nt�{q�PF��<SC��:��K�y��'[�������J�e܃/{f�$av��HHD��o���H�v|�,&�v�p{��3���F�N���,'A������܇����EE^X�?��vsw�Y ����������΀S�H3p-u��J$���4���R�SL$8��D�F�^L�-��/CR�?��+Z�Ƚ�������z�v�$R����G�>F�6יH�]�"�2ѐ��?���ٛWXz^o�.�����Ǡ;j'��Y͎3 �K��Q_� ]9�u>6�S��@~�ծX�\[� :��/��@S�1�q1TA���CgSʜщ��m%���̯������,�}���=�I�b$�.�sgP�014\
_,Nbqx�IU�B��f~�������d�7�&�F׀�}/�c���nP1Hz}3ð~�^�jI���-���(�8�K��$�+�T+
T�ޫ0�,?�-(Oz7�/_�!�f�,��]���I���2���hQi��?^ �[� ^�9��G�5��b@��e�����C��LXt��H� F1 ��tΤQ��@f�;C��#�9u�]��n"�o�쐞�Ye��� �XI�1lp�
��;IL�u�}��.x�q�_�@�n���3\���J�*l��Wڛ� �vtx�*�A@]���eo;L�9-D��I�����ވ:�a
4'$Ԉ����@�� %4�6O>e��U�]���V���9��g�������Da%�4վ�	�D