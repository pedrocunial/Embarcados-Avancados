��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c���ѢǓ2�Su���;��"d�B�,����USԻ�<LA��<@d��k�K).8�H�i��OQ�f�V�0�2.<��jI��=P�yH2	�+Y�l���b'Ҹ~��͖�(��1L�{����߀��;�%����/Wtnw�f����R��{��8ZY�? ���[zX�<���z޿|
E�zG�4��������>��3@��@f�[L���x�cPGK��0��H��=9���fz��l��}8,ėW�_e��涷py�)�H�����6QV.Ѻ�z��׿�h�7���O�sEL8��� 3���)�-�+~�ީ���uA��Wˤ4T�z�9�KA�v�k�;1��{�VP�!+0�ܴ�a�c��ߛ�f��3���j�/y��v~A�I.�y/�j��[K� �d�m��eU�Ad ��^�z���S�Ɂ58��sőd>f�(��	�nz��L<��xo�E�d<��E/��3�o{>�+Lϯg���7zs�qRJa{@-v��UWȗF��VaVBW�G�WǍ�C=h1nG؞e͇�7�N�0P����&B~��T&��o�]̤�g�6yґT*��M҆8�~:����Ɵ|!Cd8�:�#x���~�f�Lu�`C�4��;��Y]�T�"D��IIC�"K���sP- �e��j��5M����l�*B��IT_�s�Ĉ[��%�5�9����,�z/�����B����r8k���6'�������@��Xpl0���C�ì��3t����l0�rV�k�t�b��ؠ�W���=�����f�ξ����1�|�d��Q0}<Up����q?xyy�����׭�Xw8>������QFbPu��T�K�����fd�e!����8��p6]�������/�5|�����c�z�T�|�� �BȔ�]V�{
1?'�KX`��Kqk��J�`{$�/�@�����;�^����|�Ap�mOvj[I�8�`�1���J��!J��Y�� .�`���{[9�&ڡ��V����(�%_�ԙ������Nm�r�T�T�N�����wِm���u���{��a��D�j���hE>���ߍ�Ā�f�շ_�}ջ7YAh-`����?�����^���9v�8�Fr���+�t�E�?e:���+�X�γ{���A��*�y�VVs�y:Tz�a7���=��&6��ښ��g�0�D�z����:ȓ83���hk�1uK��f@G	��[�z�=w7��+�)�}��?�ص�W�/;��p�q���d��t��ֺ�(^-�v���+5<:;iƚ��L%�=
��-�z��K�x��<th]��N�q�9�`���*2{��5�~��)D<W�����*�ra��nu�q���*?oO����&���3h�K�ჵЉ"��j)a���e��q�2����N�5����y<�2�d��*l;�v�N�q�B��b3�b&�NYN_G��Pw �w���!�>:��˽
�*���wT�窮J#̴�����0>��̿N�^�
�����G���J�Z^���Ej~!��q�pT3,�c���uțP�,����L="�a�����S���,&#��8k��p��>$.~G�`��݁ϒ4�o��:������`mV����]�l��M�'٤��k%�� ;<..����rc{�a�P�06O9�ʮo�23����#!��(/��q�xn��x6۝4֮W=�ZuB�	�&�ͅH��-�c�0u?����)�@|����2��h����~���'Ѱ�~	l�տxJ�$�����O�8ĵ������IgD�-��d)��
���v��X�cfl��b1����ZV��vx�t��F{v�=� �M<��%ݔd6I$�پ!*�~2��N�GF5t����%vo_I�� !�x=j���?���<CV�g.�%�D�>��,�X�f�=Ԑ��eS;� h�A��#/��pb�$^�Isk�⠳�EkX�}U���a����t����+b*���9��ԁ;J�v_g�hsG	��sPtTU�� ��F/�.#��$.�Woz����2��M0�UVl8c��i��bW"�6
�AHqщ�ߖ=T�t|lz�m��:j�.5�ג�d���� �{���F�U9&�5,_x��rJ�f��X2�_:2��75�ړ�M��� +�c#�ub�+e�ȗ@��=��HsK�����nT���o���MV5��bOk�Av�%��x4��ymR_�o�Ȧ�|ap�`��c�ut��+{ߥ�¦�|�P�^y���ٳK�;}I�\+��4eu�,�p�|D |P3ft��n����@W��,������Y\�	ɭg�v#������G'ج`J:E�\z#�y�q�k��i����qa��}A,�؉���U [�}e��iJ~���D�������M��cDnc�X:M��O�4����Wޟ���P���\�6��k��H��7����X+�i� Y�	-��SAB��*��O��%����*�M�����[���)[���C���Ӟ�H���r�7���[Naj|�V1fy��u5�H�+iL�OiͲ_�hB�s��SBc���i���]��Ve�uOp0������-��pH7�h��I�I䁎����/�$���QT\t�B�U~\Lq촇����dg��1 �B�(M"�2��qa�Pu�����$K�Oـ(�����s O��4��s�
�b��8Ku�>4),7�*��A�%IiA�/�q�7�� �ʏ��wt����1�Dw���q7;�`0��z6E�v|r�)%�*�wra",�_Q��6����
���k���Q^�e��`�z��OvjzZ��Sb�:d]�fW�#r<sΏ��,��� Fs��D�O�Ʃk.�v�.������e|�8����֥�\�?)�NO�W����KNS'��+	l&<�2����<���Hh�2�7D��Z�V�@1�Յ6x_�(iOU�X'��⸫X,�����4��m�'�8ѵ�t�Ċx9��&�T��������[�wKQAX�e�Ș����g\<w�#�9���E�8E��s:k�L�Q�@�lb���e~�SNKd�G�PZ��k�Sn��R���e���֝:��!5�]�4�~�ahD�^�����}5ޗx�)�eXb��StW��}J?V+�������R~���*c:�'����ޞzL9P@E�
�ipV�䛩���%D�m\��Q����Pܬi��at��6!ۋ|Eƚ��b=������������(���0����B-�R�J5q(BcR#��1z}L�ԑ�r6s��	��?�:wl�r���z��7�W�� ��@�y���%�s횂(R'#����5�5^:���?��Du��.7�$,�<�K僧Ԥɬ7+� P���=�$͚U,}��M�I��A8�,L�DV�U0�r!�9F���-H✖��%�[���AI���{Q�6�ښR1&��sD�������!Î�Q�g�b�V�bWL]L������YSvZ��f�L�5�sw�$~|N�c'���?}�`���no�R��w����Tj̭���a��
�f3y��|3 ��d�����퍖�r	���QB��bQ|2�R6p��g�\9�xv��H�e��'š���,���9i}	d^��6���J���a*	��~�~/���-�r6'��Q}]q�(��zC�er�D/7���ܜeYE4ֿ`���=솽��у��J:�}^5'��6�U�=@8ܯ��:!�<�m#�8�V܆�Թid�&�-��<Hf����C;���S-�EJ(�<y^��2>e4P����6 e^SǍ��@s,��b���՟�ۊ�Ra4�o�4��Z�;�4����m�b#�.�������(���@
������8���#�Z��W3a�+�-�q�"��6w��8n���@HX�,��]8QV5���k���p�י��L��������&�Ya"�ip�%�5$G��%g�ԹS���[�W4jf���u�YIQ	s�
/9��_�Olf��`kF�h�b�M�����?�a@�i2�-c���#�u-���m��
�gm��i������<���w�P���C�"�\z�q;��!�h]�%���x�^{ �8U3�*�t��Dmu��矆����tQV���.�:>�;�"��w�I���`�����X���@��yx�	�Q�"�\�DV��\w�A�ZN\y��}��M��lUs|Z�0tY2+S��^���>B��Ad�����C;m\>�@��D�T�8`��/;.�B̰3b҅�'7�Eu�Ր0K:^��_��1�^z�&0�R�-\+��Э&x��|�����Z�7���[ϸ�`��ʖ�gk��~�k;r�;�ؼ�����Ю��V��rY�u�%�(���KE w�r`��`8!�f��ޟfD(��$b97b��*���7Od@�1ە�&}���$������|�t����C�����������~+ʊ1
wU���&�7��.JB��ĺ��B��}�@�Q�{q���%�%[y�!W+2�ّ�W��I�Z9y6 Z��� ���)o0pa�.�vx�v� ���C��W�XG�R�0_wO��սo�ʕV{�%�jS�l���Î�:��?�6W�?l���r�Qd��v�wp�k=0�&jG?a���˽8ϖ9D�y��]o��WI��@6�bZ��N���-%
�6;���%ǔ�~��{�=Ry`�s�g���{k2;�}.�����n��/���{�X�Wq�Y��m�S�^�Q.E��w��ћ��-��t�CA/�l�<�ɺ���.��9�ј�Y���U���{ ��[�@�]-�R���a-�)�	ؚ[�[�C�� ��!�(]�t� ���#�{���M�A���H���J`n�w��r�KP�g�s��4��=�,ky��uW:���V�,u��LC����,5`�/�/}��P�-���k��TM�갃��R���e���*د )�� ��Տ�.�a6�m�/���U9��W��bþ�.��)n7C7e���X������nI ���-�m����$��R %�څ\�l���H���|�.�l�}{_�*EJ�jg����Q3& ��*�R����r@��E@�5
bbp�ʻm��,�?�;��ޣ�?	V�mX�����8�u�P?K=�ˊ�u�x����#��'�</���0��ň:�	�e^';�Z���?Q��&���ʉ�j����.��&y���1T�
/�'_daVf.	`� _?��Bm�w�{���R�wO��e�������`:���$ZRN�K��uF���� �mAe��{�mK�,뢤�Q�ɫ_���Hќ�r��/�R�;�׾�����Uj�A�n����Ǉ8X���}?�5$z���@�0cC�'�8�UװT<~��d�""v�:J�&��}�G���Q�6�,��V�K�hk1ӂ�k�9�|��M�c���l���|>�7�nZq��y]4�W����e2�;����/�_^�E7-�+	@�����˿���*)��C�Y	�mۼS���x����(�@��̫���� +�V䚫ag/k�s���}GZ�;p�ٮ�,�� Xe�Xx���T���Kf�f���/|�إ�G���$S$c{52.W���n�Ȍ�4�M.�z�����Fn��:�Q��<Q<�
c���������+(q^��lD6V������*ߚ�;�j��a�Xk�z"��N�BE؊�
k�e��@-���{\�t^43߷��F"� �_*��fF��&��Dm�4����k-�m��d�H��|�6tr[k��YVn"�ĥӻҊַ�X'O~��л���J��nn~'}("�XR�#̞U|��L�7�z�`�㸱�c�D��P~���=R0�\�E�a�:˖��ތ����_&F���E�LR�_��p2+z��'�6�z�AjFj�5MB ���{rs�F|�t8������B��O���A^�N.�P���G�|N���R%.���/��+���m�bՇ��<����qh�e��*���s4֪�@,���	:`~�E�����XX"�ߟ���d�����e�ѣ ��Ջ�-��x7����^a�~��8�F��D���G���[�w��v��ٖ�cE��P;u�T{��Kx�xA���0*���8��;���*/�y��tHdzm��z&���#gaP����Qo�ܣ�uW�L���)�*�{>?���ayN��7�#�3�N�ο����Aو��^�ꛧ�W�2��:L����pq�ϝ|2����=�.�V���p�7�mԳ�m�
�g��m����oQA��Ԃ��\�h�TKI��9�V�APe#�Ъ���=."��{�=�D���q̹����sA���]v�i��#E7�`��XE[T�xcSK�O'��$��d_�]����Uf	 �k�����0w&�:<j#��F$#�j-�kZK�݊s�Y�{: ��VO�&�T�\(�g���fq�lل?3��g�"��h%)?���=�Nj�Ыٓה��{A�-��ڋ��a�:Ks����NRO�O��s;ش��;����d���{� �������/Y�L�wb��5�
����B~�oA��9��^�CWd��:�ʕ�|&c��s����s��5���G|�Ps��y��������N�/?�j#��z��Y��g��W�K4�����Ti;��ccߙߦ���5�Xc��h%i���aK��`l  ��?�2�J`v�ZBZŅk#�c�a�*4�g����#E̽"$�;,"�4�����V�I��lGS�_�x������͕4@n_F�=���M��MG<ݦ����f.����:�B�4��f>�e�Ɣ�E����  �b��,��as)!��|縘ʮ����*��3b�"�f��:�"�M��飽�n��ӣ}�<�vӞSZ_����ԕ��Ne�5���S���8M`u˔��ci�,G2�g{r�1h��W���0
���5�w�+�����i틂�!Ẁ�e\4%�B��4�َ����hZ'1g��\ =F1�u�~2\d�#5L��|��LL�X!�pp�l)u	{=���->�鞘E}-ek՗��S�I���<��{ӭ-u��Yl��	�3��Pђ�?v���D�"-3�L
�,7B?��A���@W&���߫<�v{η�.I��+<z���`YK�9����p6ݛ�Ͻ�sozIw�wX<ە��9�%ȷj�[�D0p�!� �צ}�* �\9���f��~rB��L)�F2CM�K�Ϊ	ҤVu�c��䁙F��ģ�.�ݪl��m����?4����ܵ)���o��'��D�g,�@���iuȶ�X͙�7��\ό�������go �r0�PC��@���
1�)@��-��D=h
-&Pw��~2�	�I�q�f%���A~��U]�bm��>l�U�~LݣY��.L
��&ې&�y�����K@^Ԩf`���q�Do �G�샳['ƙŉD�
�������И <�Y�1�����c�>���Ui�����a(�+�Ǆ4�`��:W�%�ޖ4g.���tݪ���3L@%C޳�,\!fG������s?���HJ����QN���k=�ɲ��TcVٶ Ǯ'8b�I������!*-Q��;���А6Cl��u�b%��u��yW6��,`R�o�T!p{K>Pt�I�u{ �s�5}1&VP/���P(P Ȃl�F
��>���p����J��3��ǽ%U��q۞���*߇o�ڥ�)"1��m)*�T����PŔ˽C�����,�m\bQ]���4�@8o�wǈk,"�&��߭~�
�X���ީ`z_�l�I�k�Z��f�����Dݗ�`���0P=& <l+�����X>_<g�9\͆lQOf5#���7�D�T���b���P��V�r���No4��0����w��H��(V�b�M�H�"��ƥ�֖���8mf��XE�ܿފ�ژH�x�9bVُ��*o���4���ž��s�����0�s�eGu�#Հ��~

��+No������TQ�=�.T�'X�=y	�C� ӫ;C�F�w}҂g+b��������,UG�~��&�2�@�얙k[	��7c���'s��J�ǧ�1�=�Q��3�Tvt:��jے�c��F �zՂG�����^nJ������E�ŀ��X���Z�P�j�I^w����w�W�­�P9o�� ����P�&��}ɡG�[��;��0��n����z�dT��'jE���i֙��db�M�m��{��{�i?ea�Cp7�0x�������O��Ɖ^ka'pz�B��E�@a
_�TP��o�^+&�,�Z�n����2t�A�8�Đ��b��O+�k���"tV�^R|�,,1�JټRu� e�_��I��n�>�F�"�m�)�����)"@N�?��z�A�֨aa�E�6�1��Fo�C���J�&MIn�>����q.k��I�w|� �b7��S8�:K�忿��e);�����A4T�%���Z٧����_w��̷����[�K:��o4ޝ���ۙ\K��%"8X�7 ^�����5�(E�^��"T�"�����g#���՜�!���}3�q��
��S>���z^��s�%��JL�Tދ2kL�J1j(!�e�����.#���7K���:��e�g��-D	.�
��̯�Rh���	��\yn%�t՚�QNN�|�@D�`]��i^\ų���0���!P{^���nP.���N?z���������B5�e��U�V.zTȎ�C�>��$ԉ,�)��nW˿�,���ŷ��a͠3�I3�B��	�f��5�tp�և+A��1�	�dQ�>�z���Iq�Ք����.�ȶ�
F%s}��pCq�3��ֺ��N�T�*ay+?Gc��^��M�
��s�����X�F�nx��ۄ��aO\���b��R��x1g'�͟?��wB�L����I��R,i|�w�m
�,|,��T\�Zj³��A�h"23�nZH���z�_�X<�"�M����o�tt���u�t���S�����=�`"V���:	ڰ�N��@�1R@���ZL�s�#K3۳���{�L�i*��.R��w�<c�^���'�T�s�Gw%{��K{g.�K����J('���V�m�l댘P�QT�e�5ݯ	{A�v~�`�C�ũ,�U|�U.�����w������^���+,5�s{�\�S�@9�A|�y���H��a�,a��^r]�֫j�M�l��sM+�s��1}p�*���Q��-rڮ>�.hϬn��e���d��{ ¯Z�VM>��x��׹w(h�G��-��R�ܪ
��t�oz��E,T'[�Jizs�W���DJ`�C/��u�h��i�
�iV)j��$q��Wb�⥾\5��b�E+x����r0�"��q3%�*�������
��QR�����a�k,0��
ONȩ����g�|1E��4�]� �e�K�x3B�'M�*
m���3��
&��jP�%�|�htL��,r`{RC��+���6��J�`��C�׊��1E������Q/6�[�KP�K?��#�%��`@Q�5g�n��<l
&�p���`�@d���P���X(�'�}��?���o��G���u�Ɔ+�&�o��S�����/�6�b�ip�d�(��`���)�����Ό�w��`q�P�͉����;�5��T~k�3�#i�����%ٻ��_Ma]^��1z�J��t9�#A������#����E�����IuPUs��)�}�~��4e%�e*V]s삎$Tl��ʰF��2<�&Zg��@����vt�L�䫰_�U�"6����E��l��y�FT�T��+�WSFq`�6O��������ϋ!؇U�MeI��i߷3A.��� �Mg��j/���[Q����SoW�*=DЬRp/��M�	x��o��"Op�o�(��7�wu��y�h��ʤ��<��hq��Uy2A� �!ߠ:ZR����fF��@+W��X�M^E	O1z�	�o(�M �\���r�	�iK7�Hz1Y?�u4}᪔h.����x����V��+��ݲad����0ٛL����� �Y�c�CAH�Fr�ٞim0c���-��(n	���'<�{�SY߂Į�G!,k[ә$����{�g�vr�F3� q�'������/�!7#b��N�<���}c�_�]R�"��׊@V6�/A"��>�\e�j�(��(���}k*��t��`��xfYD�K|���%!��8-�ӱ� Kq���/�&S���4�v��=�y���g�^�G �'�)%=��n�(�d���ele�;9�?�
� �1��#��n�\�;�G	Ŷ8�D\J�oڈЀ���g��0
�LB�-��a��S��x){�>|Iv̛{��0N�.��ֲ��XJ�dn������1��QXa�P~ >	o��n�T��Z(Ѓ_g�$�[��gr���5ک�9����?�c8�a�k��
Sw��-�
��[ԣ�h��)</�
x�u
�~����X�I�g��g �/��h�gtճs�9@-$���-5	�x9[���w~���=�$���h=�)�)�Z_�3�i9$�a�i�Yq��@���ڝ{�f
ku&{�	���_�~[]������LS�:�:u�����:�Ȼ�Y��E�!PﲤU~��q��Ć��0���42��C�gg8�*��{��C��q��'�����:�~j�@O�<��Wd�Z��ߢW�Y־]�X~��Z$r⧙!�b�>��SX]H�H��j�,�A�Ź������#n.��M�����8$?�ߍsq(���#>��~w��c���FW���Qf7P��v������]�f�V�9�/#�#�'�-���� �7�w�l�R���TY�:�N��8z���o4`$�eu6	�vb{����t�Us�JS���4�?�Q,��rp�����J4晒�9���lZ��]Hn��ك�hں�R�V�ȝh�����.ӂu��=2��P&!���O�����}��D�m(��s��7�I:�kJ%G|p)ϳW#�g;6����H�Pp�k����@)���,k������Cs�U
���F��9�~�%oζ�l�}�p�fs�y�dR����g�UN�y��׾�$�q����:R3;$�x��7�<�������du1RHO���eH�7���Ԍ&��L���P�Z�
��e���^�orzn��c��i⸑����-ҽ�5�օ�1\]��%>HKb�C/]�.V�w:Z�I����A�H��di_,ꏵ�����1��u�qx�B����1���;\�ۡ��Z_��B��Ö���܁��T=P�w�Ï���
�g�5
�D�N��Ι�=���j����Cs]���M���N@x���6����r����@�e�ݠ
�����
��8����N�g)�ˋ��e�����u�lƆG>;��:}6�^���[2�וr�U*���ӫ;L�c�A#����!�܇'s]��\�Ac{�����3j��x��E��N׽��2[���3: �L�bf�-%�۬M ����[����=��H��B��ўf��_�m�'���$�s@ ���R('��$�JK��7�4%�o�B9�!j�wauU+���q�[<Gd�)p"Oۋ�b�}�Yˊ��_�:f�YN2U�UG�)f�Gf�Z��b���Z�T��*ߴǞI��/��Rl$I���[�5
�9��@8�o��bQhp����Si����k�~+K���"| ��q�/o�i�k��`x����r�a�]'��i E6��RW?�v[�r�0Gl-�M����� ֕��N�W��Hp�d:���l�b�@��y0Hc�(_b|��=!^(���}qH,V�߼Os���G�J�A���%E_P��Ku�"џ�%��=�=��^kp��"!+���oֳB8�5Dp)Gh�� �\8�z��� w@�oqѸ�'(OXU�~�O0%�5��t��HL��m�B�&K�+�4V�"M9�������
�i%��3T������b�d�Q�Q� ��~���lWj~��9��h�a{G5f_�?��K*�Io�tO�>~f�pb�Gϫ���5#��B���2�6�T�PԦ����9���/�w����Q�4�b �l�5k7+�'��]lhQ�3H���g}�:"B��釋?ĔX���+luOw���'�Y�"I�� ���aw�[)H�]��fp~��p��Q�M������e�^�û����\U����|R�jZ#+5k�P�x�t���3;D��N"}��E�����O�δ�K��?�ڵ�-͡�|��G���z����J>%�����<?#D���U�Q1�>�y}2}LtR�	��,����_�~�*%~_C����.励/�o�Z����>l/�.�@!1�=jp�̬fE������4X�C��7�!�
ht^Ⱦ��`����58o��o���I[V�o�x[���MXQ�@��!����<7�M8oD���%;��ʳ�0Y�.��Е{)��8cZ�'7����6[�!ܫ��
��'��E?QP�>�1d~?��[LUé9�>��Žh�h⃈�˕�V�j7�A��[�^m�� �:y*l�]��� X=\i��eQ6 ���[v\z��xȹc@~����v��!���ø�QE�`P���]�2y |C��^U �7F�l%��&��˜�l3���H~���aDn���J'iށ/�,�w�*�iIE�2�{	��=)��#��ę�ٱ�N���hHIkv�P�0���a�1��1k�8���Lk��T�vN�fF��ٴ�������ޚo�wл�`I�B�U�K}&�?�g�Ѓ��� �M�K�aBG�&�`�g�W�:�� +2�|ˤO/���|����O�PQ�{�¥_�d8�`�2��B�>Q��:���t�_��yL��.�:D�{�3J`�<�
3B6)�j�,,p��=è�����Ԭ^՞��P�c[1~���Q2��H+=G��V�I	�DF����#�!��_��a��"�F]�������+�N|5��c�f	����#����L�Vo�x���O�N;h?�Q+��Kd$<}It^!^��P�=#c�*9QnPp��������q�fD+�*�x$���ȷ4E|6���r*�Fq��Y.b9��@��)�N�����4�����R�$"e�HQ�]���6XJ8�9W��*�
��,a->�~���f��Ҟ���/m�3�����f��IZ�G�W?/���A��p��)��ձ�:�j���b�CLX�7`l��K�W����u��]+��(J1���҅e����P����K>��#C�
U�ͧ6�q�$8���P>��.�7�ޚ�,k��H����9^A�=|�t�ź�������?�����vW�84Z�9��y��	����r�򠄆�_;2�yG�R7�a�������8a1���8IsBk�c�dm��6ɦ�묵6�5T�m"-#������ې����YZ�C`�D�y9Y!uDd%/��{�t�P����d�`���AT�Ԃ���.��~���7�3	�cq�� ���"4	4��]����E06(Y�hʘFd��/A%�ݞ!&^�ZYFhg'�L�)�7\����td}�����h��E�}���e$�K^ʌ��i��
0���{K����͏X�Ͻ)n(ރ�q�:?����|39Y��B�Hn7��G�c1�g��9!)`�/Z�g������i�c#��*L�b:�<�u��G۫��7�ֶ�j��Y�۪�6m��y�W4���2���T���D����]4<��O��W-� rj,!T� ��4Z�L���f�|H�&41��5=V��Nr���\/�6��3%Ϥ�9�5��	�d��1��.��4;}RA ���&�Ϝ��)�3|^�,m8 F���噌<Ԕ��*Vq�.]���	�1Uޕ���e�h�����슗3+�0�R
��_U���S�5h�H�k�ǣ�UdC�'ѫ`"+#�ʪ�%�.��GW[��*	��K��<]L��!�ȝ �a�3��pot�4�l G�ѝ�1}֖�)ǻZ�(s|��>'�L@��"w�,g#�]� ���zn�<������KB���rEleR��KrS������̬��q��1���m�r:L	��HŶjZ�ߢ4����I��ұ�խ�*��ݹ�����&(D�����%�I[�\�K���zB������JNhn+X;�/C`�L7>��U��X�:���4��l53j�
W
� �n�`�������#����;&�	�i� ��d�.}~�G$4٘���?Z��;=W"ܡ?!�Z,oXy�<#Pɓ��P�$Ł$�+�,����Ŗ�a�)��� ,u�C�u%��}l�2���'I~p�Z?}N�\��?b�\7IFdm<s@�@�2���z������: ���� @+���XW��dt�%�}b��vݷ���j伍������=
ϸ���O�P��D��F���c�ъ��Θ���� ȷ��?=��NPS[���: ![:�����9�2��Yo]�kW���t�f��gٗ��O�E ����]	h� ��mZ���F8������`��y	R�)�(��È��z��~C��V�{j�p"��B����U��l5�6-��曀,±!DY��IfɹetY���D����G��w�ٔ� ���~��g4u�2�Z�J� O~5��Y]A��&�J���t��D�?�#���%���n�,�������̞�ʍ8�?��R����C)~G���h�b��G>�J�|�ֽ"e��h��b^��`z;A*����ɅAQs9�ز�&��"��վ��RC6���=��Kʫ)Bʍ�7�r�$��/t@P����i&7�:���Kh��ʼ�:���So&'���U[�| !6B��� "v���r�g������PFZ&I�]�/�:�@�/�F��i[WW���#sͳ4�^�w�gaMw#��"*����i�����5܀=x=�el��7�v�8k.�-�_�v{��6������w�tB�-M*���%�y����4q�eKk�����$a?�4�<����e�Yp��Uռ���S�����#��ΪM./�����o�����T֦S�W/��C��u��I�Hx�I�/ތOԤd1�c�H,���C-C����z��j�a��u�i�*����1W����G%Đ ����)5�`��a���L���~��L��7�l�hcn�4�N�Inv1vNU�d��k�%q,�`w�}��l���VˇC�6 RO��s�G��sHfĮ)c��rȎ��&/�AU��O'�\f�t^d���nM��<�p�ڒ K�.�2\:ߢ���Yp���H��ߨ�(o<⌤7lY#�{R�[@����C�|��%������z|#=���$�=n��/��]�HU:ӿ�x`+_���־��/a-1؏O\R"|˛>U�!�%����{`�$�i)�qn��$L|J!L����O�9!��)�N��9"�8u:j����� C�6T	@��R^��T� �:),��H5x��B&�k�W`K4�	Ь������L~M ���R:yH�z���%Ѡ!m����9r��<�PX�1�rB&���W���DSS]��,M��܆r#	��џ�ٔ�mT/1� ������>��۪i�e��Q�=�R.�>\�����~)�����`|m���7�?��m*/��S5��*�W{o�D�mLĳ�G ��֫3�>u�*��ǎQl	�j[�=����'����/?�0\�o*�,�z� ��l�/#��a�.� 2;�$�F�2�`��b���?���Y`+F����tS���B������M C�w���^��:\U��S�By��s�&͵Xt���]��	lX����R�j*�]&�����qr��v���w��/�O�G6ԿY!���Wę��@������ ��?��|��	A��S�X�$[[��x�sŮ6�X�A�b�l�@B�\?l���i��_�	�-o�7��A�ȟ��w�`��*MG�̪��4�m�GP�we<����%�%J(���|i%�R@���\���;�1]E���/r�#���������IV�V��#���-��8!�T�UM�T[�{�^��3񬖒�⟑h&-l���G�	Gw�R,F&x�])�8��{3�)�j�ɰ�Ǜ����~Տi�9~|!"��*�X�.DA�>���7ى����_�F�����)9�꓀Y�;�]��V}��`��i�0��b���@c͞��`�S��\}��\���<�Q�g]���k)０�u��K�U<�"]�=Uʨ�?�?���^�<Q�'ː�Ϫ�*M�*i�$!�$̜m{�m��r��چd���6'bV�KE�ǹ�O�ޛ�����2B~���J�)p�n��$�#,��#�?��A#c]�ߛ/q��q�8豆��G{C���Rwh��/�b)i�K
է�ʒL���e��gb ����D9N+�*@��)��@[�����Ō�-��"��L�V��sV�ԠiC/>N�A$�x2S�G����|�e�1��}谛��_����0p9���B�닿���Z�o�(B��Ͼ`-�1�[a��Pfq�QX��cF�9�*�F�k�Y��M�Ʋ�F��[�BQ��3"��a8��D�0�8P��䀓�⦵���#�a�ځ�6�;8kEt��װ�����&{��ڴ�vw��,nP���櫽�@:=t�'"
������l�fx|Z!�O`L��6�|!>��:r�sI������.�m�T�)�&��Jv����/�T��o�)B$(����k���v��6X|�dj�Q�����8/���p\���ʗۮS�m.��x�I9��Ƈ�s�q�sq� �5C#,1�������
���NQz#@�C� �h�W�抸2�7�$��8���-��ڇ @�Cû�Єu6��px���o�����5�S�X�R&fO6�Τ���Y��=k&WTD��6s�Z�^��nw~e�0��e�!��ˈ'`U�PK
46�-A��.wI��;k_��r�s�<��.�y%1��_�@�nz��mr
'	�?@rt�g�Ǖ�s�� RMiCv��#%�8��o<i&*4�STf�a�� �pYs�å�r�7�2�W3�0G=,P��#���i�a'�&�|!n�ai��-�b�8d�Na�����I��Ӈ�Y���m��Ú�_j��"Q�{i����A�\N�kd��V����t��+澘��<nU4c�U��0?%6�nI�휍���^ �A
�vK��jP�Խ�紼�=&�N^�T�+����&j�#T��y�ɬ��V¾����1����d(������	𼵨�<U�N-2�&r��O�p�ޮg�������ì���7���£_B*�5uȡ&�
5�O�f�z�F����{��"���^48e�0�A!z��N����l2�`�ZE14��*OL�$|P6��-�A�)���R�.u�9���H��F���b?�S�Ǆڡh�Y�ff+	���6HV�:�?஍��U�}�)�G�{��>�nñ�j.�I��yȀ�f ��֦����(�Ev��&�;rLAa��M��6Kw�&���h�\��v1W������md@�(D�CC�<�4	q�
Yvm���<��k_�36����F>�[�=�/��4哭�APu�%����XĂ�앶vA���D7�Sp#bl>�a��U-ď�K&ǹiZ�����E}�R�>��q��r��D���������)d4�gx�I�@�I�^�?aA��l�a�fW�?f-m�N}�����;��`J{�|�&uVi�;@��{���L>�\�ǩ{��Ek�:�<�	qy:�x�h:�P�l��#A��p&'53�F@�.�o���\�����FR��0���&��5�\����(^��G�-S���]����X%��?6f]��)�( ��Ћ�dsЃ�%Y_()jו|�b�Q�k#�����!�P��߹�Ŕ|R���2g.q��L����96<�g]Up�4p�,z�i^�1N�%U��ʋ��x5p�:�L���{���8��o�r��T�@jx��(_���%�F--ϸ~�������<�'	�&�WJ���v�%:�#����!�n�slN�>9A��`wEPXl�m`�~)�a�V�p�����/�����ы�gRd���Ce�z�|�:��3O1�93^@ ������9�؁{	�>�H�/���FM���ج��$�i�ٽ�Ydg�ţ@݌���:�q0>���&�4��7��C���h�_�v�������;y�-�|�R-�ᱫa�-�:�N�F�z$��f�뉜Ѳ����A�����}|��3�"O�UOG��qҞ�Z���U�.���Co����p�]#c��@Z#�Y��?��j�ڀ�������L�Cu���G�5�USgx"�eX��N�߾N�7���O������fZ�,Ӥ�P�f����t�|���\( .�S��~�f���wW��f��$f���{�sKR'�˿1"|��B�zl���p0����*�7H��&ݭѴ_#����'�8��v֠��%��K
B��8�\���݃-���1A�G���vm)4p� �l���~b�4�i�ͷOa�D��}��Dd�1���c��Po�.S��*k�V5�*��H�0��Kx��F/��N��_��G�eFcG��OE�ɨQ=�BŴ�n��Q���z��JAr�����?�ݛ!;1�":ƺ\%�ˑ�}p��r�̓��4m �z�}��Ρ��Zԧ`���o�i�p@���w�Lm.A��}�ڷtgzS�s�+0CR�O��oD�C����d�a��%F�$"�,	i;\�jQv�F<`�K���AK�7B.a��u���N�(Z9�$Um�!TR~�@m�m�d�I6��+'�?��'f��s���A�k�U��Ne|(�Q��ӊ���Z��׈�\�ݴ��QK`A�V�l*/I��c����V����g=TͿ���r�@��Y2��yr���~��i.lX�l�~eI6чc���r8�xC��V��Oϴ7a�r���6Z�'���h7ɳ5z>�`�8��m_'��7�>%�XNj�w!�x���� 3�u�5�rg~�M�K�h�Y��pŨ߉_�J���E��:�O�د}Ҫ��M];{�\T��4mL����k2S�Ft��B�v�8��lSJl�F��<�|k�u2����ҼZ�nx��;�ƨ��_�}%}��>��t%F@/��^b�j^,����2�Ȃ���&��_g�j ���p����߭@�\���S�"�;x���~J;δ�֋�õ Z�J���ce�Ňc!/�8G)vV�JMh a�I�����q�+��:�)E1����-�!�oCR��rc�hpT;Ċ�<��J7����pz����	QѾ�k�6�2t[�A�������-j�h�Q�X�7Vj���Ҷ��:B��fZo3�"P�����.bؔϫ���)�T�l@�q���g8��S�>�{�^���{#�1�,�2�H|�S},�����`1�<ґ��%�-έ��V��6�r�����f�y�~$R�B�Z�z1'�`RF�u��1��S�}R��0O��=�]S��nB��+W��%�:�mT�up5�]��֙�OrD*�c�Z#�&�'lu���!tV��̗e���^��/P`S�s�hoM���IZ�W�0:#���wX*A��D�×NEKcF���V����X�Klˇa�1-�ϊ ��Q N�QZ):0�M.Êt�QuG ��if�OtAۇCP�t���G͌?��U���/��1��E!Ъ��a�KS>�o�H���&*fhi�7�H��+�8�W_�����i����H�"�UBN����FW�����B����*�P1F�>%�Z�	-��k!	���˖I�\x�����= ���_̒��IA�|�a��=St,�NM�S�WA��SH��aq�I"Ғi��{I%F�fдn�Х��?i�+X2(C�X��@͐�g���Rvni6�^�}8TU����������&�xe<X��<sA��6��؎�u|H���8��}�QJP^�]
�H��Z��^Hf����ɂ�����-����3�.;�N�y֐�y�	���/�_ֶ�*ռ����e�G�4��{�3Z"H�=�@�ϒ%��>rSԜ̐��p�t������~���#��/�Kɷ(���w����F���a�t(類�����Q����-{��}���yϋމA�+"��F�N%��ɴC��N�mLH�r����=~��?Y�
��a�,���;yΠ��vsҗ��2:���A���o^{~��*	
��n�h5[:)���[J�f�����W��볥�j��m� M��;a,6�W#�۹�P��Jr�u�*u=��{���FR=\��)Fɤ�V�����=�:�6��=.�+�Tl�߭��l�h�u�y��@�қ#�!w��0��_` ݂�������cO5vd2�R2խw�w�M5�Q%=�q�/�A4�b��)����b�fK�3x��=8 �y�fK�ie��^��+��z�33e�4�H��VX��b��
H��@o��'`��@A�W�a3>����ʈ��K�$S�4�F�/��?�)v]ύ,ܻ��"��D��+�HS~�,\��4l�9��,3����4��o�"�B��rάټH��PW��3�o�k<J�݊>⿥���
���Cm|26�=C�͋5��/���)nP�3ݹ�@G�"�2��C4|����m�N��n�8pn̗���c������C;ؕ(�j�f�q��A��̵�8Z6����m�$�/Ȯ?�ٿ�p��DB�/�3e�V�7'}�~_~�<���P���1`B�~ i��M�o���(���l�-�2�&ğ1;+Se�p�P����� ��l���p3��G�/r�)�|�S��؄����7�u*�"vzU��ye4��IBTS�X̭2�[>�Q2)�ZI��?Q�&�$(��N�X11��%�����������9��u��2�y���CȆ#�"@�n�]=:�hR�@��.<�ű���Mj@ɳ����'���(�`х>�ǈ������5{����N�>�- n�Ô�F��7���9�,xh0��ት�p�HX�D���8��ŝ<��,!��^czU3��|�(ty������.i#�{`OQ"0��k٠��k��-:\h�v4� �ؗ_F��(3_Xn42�{�<}�L�#�ň؄>Hbҝ���z#��$�2L��S�N�I�q_�&����3�)@��XɪP��IH4b�g�bh��Q}��kB�8l�
���&�:F6�@��gN�EXU [�v���P�CY\A�A�	�)�����Wr��]CL��|����&x�:�����ޔ�*JNeΫc���ro��M)2��k܈�n�����Nnf�;A��[�H8�.�]�z@`��5�.��wz��.jaʺ�mP�΀�Ʒ��;�P��N�*\o�#��ф8�η��%q�=Io�}&ٿ�2�)�hPté�c.$�b�V)LN��e��<�*f��v��&j�Q�U4��>wK�P�y��'����c�r@�K9����-�V�<"#� m��u�zz��N���M �)�w?ִ����Ź<6^���5(�bTg�T5I�-�G1F����8�^���MQ:S
a�hEy���>;�>�OD0@L3�+���Y(ƅ��A�w��g�0��Khf��V[�2%�'���C5�������mvoӻqŭ�;�����j_��aiG���6W����P��m:�K@�h�����c��kI�9�ֈl�ێM'\aU},>f<����2�_ߗ�[Vu�v/ˏŶlݚ� rY~�|x;������2p\���b��y���OH� �I-�v�l#W�C�4m�Í%�T�K"A���{#�Ѫ#�\-���Ff��dѤ��� �,������I��f�A,�f�l�yE��I�6uk��!�I���P$o�����Qc�h��h�)f����hnh".2 ����ߟ$��!�#7�Ef���������̩��R�3}є_`Y�>��1�r%��5`�d�d.�x�:���F�o'A�;�]�Pã'!1�2g��� �BD$��p�W�y��;�N4D�5��W0`��R������}!��e:/Һ#7V![]��,�Tb�ʡ�]9@�GT���/lN���(S:�`D*�R�=�h��U��ImE�WD��\HG�����i�C�ε��D�>o$�v��� F�[�s��iR�E/�)���1��ze���^E��'Mr$�atp��ژy����ٴ�8q@̔�n|�&��;/�5�(��D0x G��mp<�ܔ�(`}�YOb�[�8����c�G��?T�]��a����'O���e���EQ�M��.u���WHˬ9=����:	�1J;�?U�<�|�qw)|ke	��{���Ԅk��OV�.�~<�]�tT�:\B���O+�H��D����k���YzX�%-�u��_�'j�@�	�b�^-~��d(��b���L*n�~O���&��r,�g�iE�|����m������j.��X���f\����?,���N:�X�0]�!���5K��,gQ��~'U�R�^0���xf|�RPS�>e�c�懰�0��ʣ��L/���t{��w{�{�`�yA]���4�F�K����ɜ��UW:��4��OD�H��Qy	&)��4(��л�PK��2Qw������j�]���9��\O"09�h�G�%��B �['ʢ�K?�|�G�>��Q��z�s�G�
_����Y�q�Kx�r��b[/�)I��o�&�w|k�g���k��zH!����"�P�;��K�&��2����(b U?x
�H�~���\��:�T�gn�0D�J�`ݤg3PrX�d��6��͌X耧8}�dsj�x���(�܉�Un9��t}ڟ�=������w0qP�����ˁ	�Km=P��9Q9s�%�F�E��d̘%�����u�"�G[,�1ikJ�RQÖ�Y���
���	WW��]�������D�z��[�z|��2����p;"�y쯦�>7,J����%�)�g��s�ZS�b�i��������������j�<�7�bݬ��/��chd͍2(b������q��� ���6�T�`g��_����$�f*�$/pL�i���S:�rS��K�� ґԯ���2HE��	�h濴�wt�#��;]�p�2������VR�Q�(?��0t��1�0��eẻ����e�oAISp��*Pg;��V�e�5���bk�E�+`����Ҁ))	}��9�K����N��2d�i��VV�"O���d0r���b�Lc�� �n�F�Sx��NZ L�E�=Z�t:�{��&�
��aW�\�U��٪���	x�i��K4�#2wl���<��/@v��N]�����!I�H������N	�£z=�� �w����U�����<�Q�m���Y�7.��+�Pv#�5��u�C���] -T+�$��^W���	zS�?=�=6_�^Q-��,;�O}��5"�;���_����2�s��>g A$��1����rE����i�WS�=p��I��:���<���#����ǅS�v3��"��o�@e���&U����[���V�~=f!��k�=��*�Oɶ��KP$\��P*��[���_]Z|��U�L�v{�3Q*���0�ژV�����H:lFQ�K�1�0��,�V��cH9j]V @g�̉��SM������y��6��#�Rx��2�J�ME!m�DH�~T
q@����Vw�
����I��`.�"�|�%�kd��|�,��B�h�Q�έ�c=V��5!a8�㋪�N��Uz�ֿ.@
��;���������g���i��d �J괉�2�Eߝ�:�T%�|��R�̯����l+ݬ�(م�V
w�FpO�kK�Y�O������T���L���tQ���K�-DŮT<�h4�F!�.VVk&�+	���/+w���E�L�P�\NF��él�am�ķ`l-8�~�����`9��bZ�0�����m|���:���� B���}�G
����Z`-=שL^�(_=�I�0[lT��DR��8�C�eݯRW�B2݈bTM)�7�q��@� 1Ik!���oH��jƒ#nh!�E�G��m�Am��1�QL'��d�@4�5���n�aCI�*�P��(�d��m�(���v��V���Ֆ�dѓC��~����͵�E#���b,�f}�5�@:z�� -	څP�q]:1=|�_ݛ��)�g^������.���n ���ژ�G8��:&�Y�5 _�����F^wߺf��r�X���C!{tv��w��$/�Q���"i�Օ��^�qw0�w����>V�6�&%�`�Oz����2׋"O��5*��_�LNׂҲ�ʗ����$��~�[�ڒ�j~e��`{���'���zW��7QV�M}�y��-����Atp�2�D0hr���E7�(��HKI�xC���C̚���3��}��W�5�UltIi����D��	�����!��F�2�th��-(&��cmb�rQ�S������rV�U_::'��30]�*Ӭ���	7z���
݂	*���$���F�P@C�?T5	a6��A�ʪI^[u����X����Do�x�\o�X�qG\zv�ըKT�;�b�	�e�`��	���HM��c��D�[EÒ$�@<;Anf����릜~G¹�5ٷ��j�v�a8ړ]����U��F�Ȉ�;��'rm)� �=_^@�%�jʼF=��@g�wnJMb���]x�7���|��|j t�L/���⦸j[��'��'��NvČ�������S�^u�+�$���Ւ�ѵ���K��M��hN��x"��~�nV��F,��7�:-�]Xp��g0�U�μIcz`�N�,jt��6�S�Z�0Ҕq6:�K�!��O�$l�]��hf�ݐ[22M�LkS�XL6!_{r&�v\�N����玝	���.;F{Ci��;�_�C�5�;M�4u3l�̋	�t�عV
�uַ�\��(��7��2#y*/P�m���&|��fq۴���s�rے���uZ! A��j��Ꙣ�qu��bWT���8���_i��T!���l��0ơ���<�%oRXw���hߜ�B�#U����Ux.o?oG��
)s��C5!�х���6�Ot�6���9���
E��r�݆NM6��[��E��ݥ{�/|�P���7a`
�S�m�sNx�l�	z�i�4uc�ts�T0X7�F�K�l@�*�{J������Gr���+�p6LX�nӰr��ICQ�O��U��f�e��f���`S�<�`�==2��Ě ��`t�k�VXY�.������+_{|��O��bKh!$���Uӡ�Mh)�"�ꢢrrv�i�� �I5� �*���d����xx���Ԕ���wjO�����j��n��%�
RN[���0��R���D1F���Z6���^���V��[5�?(���*��ޅY
�s@L4?}`=�3�ϦLK\wcT����o�)�te@�q�_E1/1�-zQ��	G?�C����~F=5��ࢤ�1Y��I��f��>?��?&t!�}Bz��q5}�-٘��z*U�kԠ�
�o��RxC�R��E��v�-��2��}ЋD�[�s� �d7��#��Q�3v���Վk�H�?�T߷�EA�2;"	�_��Ȱ�Dfأj��1���|O��l�i�T��P�@�qwa>7���>���*<��;�u���-K��E6ٌ,��g�֕��~���<�p��duj��܇og���A�/��D�d�q_�|F��s�r�����J�f�xZA����:��z�ׇ0ԽBζy��':�:�J��e�M���	��p0�,_0��N���_�:����&���ĉ˜g8oZ$���􊆬��*d�i(���<�f��b�<B�r�a%��=V!�ʙ+pK*���a���$�'��mI��nD!D�����J�DQ�n�F>�ǁlO�A��W>��5/���0��կ���y`�z���:��X�N"���oG��'3f{���Rh(�ͼ�;'|3��.�j�댘�ȼ��I�	�d���"�}Q����W"��<^�O̃�����u5r�9�N��������|�x�(g)�N'�+J���Z���Բ>���J�j{�دĸ�c���Uz��2L�*����!o��ś&�1*�f�-�]$�瞙
�[k�&S���
(� ��O��+"�TB^C��J�@��fL�m�Ă�X�� >@K5�g�W)�}���w�brW騚�r�߽d��;�x*�Ǎ\H渷x�E�.(H�5�-MIe������g�[Q��)��ޠ08>e_t�a��w�n3�H1a����Xo��X}�vv�͕z�M��
't��y���9a���#w��χ��Ȍ��8۪$�̣�n�锎�S�MY�g�U���R��20��F}�%�ٞ'�
)�LZڣ)~,��nK�([{�MN��fX��7��9��U�]S��e�3�Xj�`�1�ʺ�a��t��`t:w�r�DM ��z��ȿ' 1��˜r�4 G���Zx?��v�Y,����)�ev9�3� रO��'Ύ���K�X��W5,�NGq�$8��7K���;C�<?�;i��6}���:(L=�{.��B����M��;���6R��* (�|�� Y�7�z�_O C�W���Bb*��Q]����3�my`�B���&>�I�Ƿ&�a,?u4j�3F�4;���Bm�sV7NB�����K33����&`V3��@8I!�-+��9���S�DJ5�	��9��U'���y ��EK�y:������`��byPlJS5��K���MD���a�[7�!�І���>G���:F�!|;=<��6K39"r���5̓��� �p���H�ezB.M�� �h���_a��I��ޱ#����L��3����Ũ� �����?�g|+`�?������'�8��P����xq�߅�R�#�*;�i�9���:�A�E�P(6�O��'c�͍��!X=�X�b)5zB�ٵ�Tŉh��t��Ѥ���f��C�}�A���e�
#�e=k��T�C踮)�5]�<�&Y"�{
������dr�SVd��zF�e���nO�������b��Ğ"w�H��s[�9��D�����MV�.s�?���Y�	BG����������9K�o�e���8�$���J�"e;�a}�G"l4���(茕�\����ޓ;x��J�<R�o ?�����Y"_�H4$Y���U��'�>z��+�tg�s'7�����)
P~d|����u.�����T�ۀ�U}Q8��kF�;g��m!�\���jY6f:cH ���M{�}���-g��R���Ј������A�QhȠ��b[./G�2$��� D9*�G?~��*��.��[׎ߋ�1.�[�&uVk�^���쒟V�N[���^�Έ��m��#���Cc�q�rd޵�t;I`�	lz��b��#�T�n �=ّ�ײޫ�oR�d{���e�A)I	۔W�$�u�� �{�n��I����q���'^Aa����'ޏ/\S!N�#ˠɵ�G��<q�{ ZJv1 z�6�ּ�
4�>H�w���WaBP#N����Ŗ�e��-�^��YM�Cɂ�����9���üzȣ��R�����l'4�0o�
������^%��B�|)��)xuu�wL�J���~3�ʓv����IQS�#_��1I����쿃wE,���Fݽ���w�Q��g\�y�����QMR���h߮�/�O�]|ѻ譒��A9�9m-�� g��k�� �EFf����U��+m�nC,p�ؗTp#b�N��n�u�QN���E-m����ß�p��03��"��q\J��-�$Jч|)�ϓ�3�$fK�\�z��_ٍ�\0�x��~�[��9E�;��e��7�.)��Z���ig'f<�/Ƭ�1�	��T�$F˻�x�k���p��Hy%?ϡcN��Y������d�Q^��G�&=_[�]g�V�h�o𣜤4~�b���讛��5WsaOV���y O�7gm{dT�W�ZL� �_~Ho8�T�&�`�NY���-Q�tJ6�B�9d�(��Z�s�H0��jb�Ak�N��ތ0(�QE���y�Y�J�E��TK��[���L"��]���uJLF]�-�$﹀��,F�1�Z��#�PL[_� ���n�uNE�K����	MM��t6�L�yCi�&_��ع��b�up�S�� ���u��>��iA"!��R��@ȴ�n��d9����L#ÁҊ�V1��Ee��>�~��� (�MaԱ *�8�XG�G���������7��o�z�4'2��8�յ<a\�Z���4l�F�sH�Z�=��r`U��㫟��P*��|���Ǫ��̌��(R�� ��,��Q�vAEM""�߆�.�`zg�%�a���t{zoV�u�2g�}3��S��V��S�I%���%�m@F�R�<<6�����L��ylv���%��Vrs\j�9:h�aC:r�`��An~��|e#�N\�.�8���%Llϙ����,yT�k"L���0�	�2{���r�H�ھ}�F� �Rt훧a��T�IKo�X��"��k�i𳹹��2+[��@�a�P�c�̫���r&X(	.��Z�L��[ee=����5�?2����*˻�d��ߪ!�X�|�u����Ke5/��7Ο��'~w�@�A%�n��#-{:+<�+�����meJ�� C��w��C������+�l#�r�!���1�v0������n�}+�$�w����k)�~�.8i���:@"
�G���s�j골TgZf
ŉ�߄�ި��[i�'��L�׏
�p]5�*���L�8=��Dj��).��>��x�0Y0�ϼ���%��N�A�� �ޖ!*�*����i�u�����1��zQ�&Qcc���o1��DW
xh��%���.���:X3�l�M���lc�i�
���Q������k,�TR��Be�F�e���{KH��^�	,�����I�*S�T�w��]�Zz���wG�r=�m7J��/��Z9s�X\�(2�oJ��(8�(�ri�z������>��p]<�?wh	>=�� Lb5�~^
S����5�X��u�P-
��;�~��1ǽ-N�b@�>��*c���=�A��Tr�>!��Z��+��b������N�+���T��1# �ƻ-�(�B/�P#���q���> *
�&[FW�<�%��U+�^L=qG�v�a�o�h�zN�ɸ�}��� ӟ�tv��Ӑ�S���6�����������L�B+]�����#�?�DuG[s&�D�U�6VV���l���V���m�]�����|��R����0����HK��S91�\���(�oz�=�P]sF;~}������c��'>3۾�s^�.�&w�˙�k!*1�ڹ;��������5���_���j'*d�a|)ȕ�m��Qi�P.���x����|��:���y�o�7�_f.I�KC�~��I����E�����vR��1YFw�w�$	�q���)$s�n�������	�@јP-#�����@�Ha���pUl(�[�nǈv��M4�^�2���ۗ-`��.�I��v��Ld���x�=W���Н���&�.�qc���d:c������Y� \4t�#)��Y��z���qսyJ%c�C�6L��X㣅���Z���;I��n�ƻ��<?x��1Uq�Sl3��cSJLU�y�� b*�컦J+���G��%���.�����3��aӣ��}��yz��pz"���!�ܶ��C�A6�Nr���ߜ�iYS���3U��5{rm�:H^V�������V᳥���0<
����D��p:�9��K<�K]��ص�z�J���Sw��|it��RL��{��A��I =S��g�.�)����7��g~BN@��I����v^<0�=�b��a\���I�9�ى?�g菤#�ljc=�Q�'��ʧW�o��'Bh�DX�f:�%$ug'ö�Ȋ����.�/ђ��N��:�h\��O����*+Ei��]yɭ���Q�����H)|���w'K�<�v1ьfx�l�U�S�[D4����ץ2طR/� x/����_���:�0W�
�~F���S�Tr?����:��h������jSNlX�� e4�6�H\!�15��ɽ�eW�I'=!���v[#lj5��(�δ�l����W��G�^:�|�9�p^~����� �b.n�_�a\C��BS�pk)DBLV�l�-� �Y���M憰�1�,��)z"|��Y�%��S(8W]n7v���Ƥ�L���?V"�-,���F]\�aL֢AOJ&R|(��7پ��w�������=&��)c�q��?u�+u�/�y8�p���0We�)�bW�7�]=����)�4��`�ϓ�;dP�v��Z��Z�N�M�/���lt0����hθH�Ctɟ�h�3}���{��W� r$�G�w$��]%^}zw1
ir�����E2�#���"k ��H$c��<��M�n@�zH?����X��8��i�Y	�:�F���Zj����$V	���c�bB&�_&���I�q]`��RHl%�,����[L�h��F�U��g�[���������c݇'��H�z�sl�ܼ�����#픊����麚�+�s�����vS	��Yf�c�~��M�-��RN�|�c�Aw����^"�QeY"�OQ��|��~j��Z���)���@n�r���C���Q*��Kss��>�T���_�7�� � ��F6�{�q�����d(� �dŶBU�/�e�������
\K����-�Jf3���p�tز�5�3w��"�v$
�[Q^��E�)�)q����Eft�OLq��ʨ	�����I���/p��Hp�$T`��t�q��
߽n�O�G����a�"߫�9.fK�b��xq�ǯ���L[�}�닖�������Ͼi�Pp�"�hU+B�?����,J�8� ��/�CE�?�Pk�$�>��,�{
�~f��Ľ�uT�೼?Y�ङ�<����|�Z�VR��`��j���6{�K��Fg�TBR!8����Tx�z��G1��d�w�<��wW��c~����#gfc����+ZE�o���¦�I��L��%�u}кm/��`,+�2�(�ܤ���Գ
���T�c�nANX]�ri����C栂a��k9�SE}��⛨�Ŕ�B���]���E�9���Z��6�@��e [��k�r� ��*��s��?) ��E!�<4kh��[A��:����q�¤�KJR�j8}��X7���F���8�B(a�����<��Vbv��?������q|�
%��P}�8T�<[���a���M��o���:�ݰ���\�0Q��U`��
�$�E��.�k�?G��Rj/o�1�R��iY&�]�r\ON|D���nٗb<[�TF��Wl֗�+��/�{��'���YT0��k1�����j`G�j3�,1�����[4�S,Ξ�a�7���;\p��V�Yٓ��N?UWWQH�3�T�������G���gH]D~��|�z�P��aڒ��#�h�׌n�m�'~�!�1ֽ�2�i����S;�,c�|u}3������u�v�a3|H,i���[��)������ɟU��(���(�� ��a�c���=��J��}8Wo�ծ�Q�&�2)�#���e�μN�j�B1���l�i�ϛ���w����ܧV5����a�`pOG���,�u�R��(>��D�?����$�H�!�^SV��&uz���x�®��d-����/H�ůef3���)mb&�[*�s�f�L���D��x�6��<�)�<��$�����h<$���/����e]|B,Nd������EP�h�r�!� C9yOd�{�~P�l��E^��C|��pڀcy�����\�8&�v��>�95�pn�*��f'!@zvJk���bimo#�[�\�L.&��#�Ƨ��2w��Y�m�4$kn~sD{���b,X:hk���"���H(��~d�L�!��&'����j�Ұ;;����R�0��M�}W߶]���K�
��J�I?S[!\�^�>��e�y�Fi��}���OH���*������� yߍ���eTw����):A�7r��zZz&D����h��ĝ��|K$NU��D)s��A��6��ϻ�Uz�&�m�N5�5g%�j/��Mi��TY\��v�(��<�*�؀���v�Xlm{=�ɬ ��IƁq��o��v/m�տ�3�X��l��+�'oB�!(k�H��f�C�����{n�3#
T�s���¤�<��8e�տ�F�%1�Jx1LCi���R�9�c���m��"S0���	��Vf���q�yE/�k��͚C!���j�h0���������cֽ�g{����v�#������}�Z/�5�H���ls��u�{ռ<j���X�q�~*�}��>���������[jП 0�\,>����GP�oҮ3���8��QT!Kռ�:y����D���.np.Ł��#�
��B}v��e7��(R����������ީg0��I��h6-�[���̧��>���v���}���*�Ā2{�p�TT�6Q�<�%a��^�S��#E��2TKl�y�&�H
�K+�Fa(ٺ.1n�Ët�Hcs�*<�n�5�8��8�_�<8}tk%��Rk?[k�]��W�j����ۂ���v(x�!6Q��
Q���,�#��qJ|
w1un`j�hQ�Y��|�JTO�A��*ݳ������k�5G%|�7mú�'�dh���j$���i�d(���b�ܙ�i�=��i�]x4R��\f>�Y��E�R6$��{�5.�h8���%�]�.�.�0V�9l�鍶$���]���@��8���{O�Fq��x�J�`of��n&�̻�\C�p4���5�RB�E�f�:w��Ho=�����]��D	�泔獷@&����[��IY�Y�owN�	����ń�o�����?��Kc�)���T� �b�8��f�6�+ �]� 5���/JF���rInW�	��<���l釡����sU{�Tk�U����'&������S`�b]��\,6��Y�����U�)��#�;����W��BgtD�bX�t��u(љO+r�@+���Ԭ��`e;ƫ.i�ke_�E�����1u��5'���h
׾̡W�z�p�߫ğ��-Q��Nθ�k��h�s�B�ɽ�v�2�ΫOy��T��AF���!�O����Ͷ$�ޥ7��%I�B����a��� �I����n�<j�����S�A}��)��<54�6VjCj+����je�\}M
�bg-�ɽ�����
��NMa��0�S6�L�A�n�(.�D�F�rk��j*��e�j�s�?����pk�.f���Hs���qv��P̒xb%p?��9 ӫDb�A	�%n��ɼf��L&�fi�Ԁ�u�� �g���:̬g�����B�z��k�i�}Ԩ�����gf:9V�]��N.yEN��n�����/��?/&d�6u������A���@�d����nHЇM{�w���;�XC\�8(0e�T���ь�u䧋Y�+�]�� ui�lK��u�s0m���-�~:��a,��#�/��<~ԗ�6�4�K:��dpe���*Lo����N�} ��
>@���c2�t�\E��^����/`�snMH����D=�Xt9��5��m�,M-F�"_t�r)�I?���q�H�F:0mz}ֈt���!{y"ge@�P�U}�ɛ��j �J��d 8��dl�TqN���e�����w{���c�-���^nR�C�{|c�u���n�E�a�˛��B�^�ͤpl���=_��=����Hϕrz�e�1Q�}��w�u�̸};Rf��CV������HwC������"pH�%&L��=ع�g� ���'���,!"��N�&�����ez�"�8 7�������m�q�Aoc�u��:I�?I^M �&����p�oD��&�2\��߉M^��=����M�V/V�@��|�D^'�3m��PA���v��5� ���EL�+��Է+!�,HE93��~Y�W8*�m�(\�6)/	��2��J�z}�:��a6�	O2P+�F�1mK��upe�ѕ���P��W��B��򹤓9hU��^�+��ΘS�#��>l��Hp�ͱ��I?l��'ģ��Δ��-!�A�J�3Z�l������*�X�e��h㌟~z@��^�V��h��<p7A��Ue0�dh�Cߺ��J3�����#9}�X�3�kP�6�����m�������:�js��ˊ�@\�-~*�,|1х*�ZҖ�dx��Y���rS��w6�y{MX��s+\�޵h�	��%����V���n���l_k�%�@��L+fyu�	Sм.'A3���|��5\���yn��i%Ao���U�j�j�(-���~��/eޓN�줥)�:��v��UM��+�^�' 속VR}�@����"�cR�>���.�ʄ�p�=nBv���$P��h�&+^��+����gL���0]��.��HZHa䯀޸�����70�x�PŷCc)�LX^�ș�9�����o��B�K08�3PEN�T���d%���ԗ׿/�\���l�0�x@f�Z:]ϵV��K=^��Ө�^�מn�%��ƨ����'�>vy�!�j�:�!9
������6�"��Oc<�n5���z'q�#����-0H5�Ћ�냆��G�z�K�M���t��Y�p�,��v���<�)8�⠂#NLΘ�c����|{R�ץ�X�����L�7WN/0�(�𤇡���o�������	4�w�G|6�������f����Oqf��<.�$��1�yq|�Fx�� &c� <DJ��mX�no��B?�-qR�L�� ��J&�޵(��*S?FT����_V���A̿R�l�?��Or������y���+���)؟A���R��}�io�:��U ���}�6�`��C�~�rD��L̽�.ͭ"z�a����?p?n��t{oI�&��ΑT�����'�u4�Ns�j��@ݫ���C�(���F���2|4Xx�.ڳy�79�n]۸%�L~[��~��i�RfnCܑ۟��p-''�#��\t&��	M�T��1��[��X]���2Dv������&���&��ʈ=Iˁ�'��{G��1-y��.:1G�T�7-��������
��P�ݿJo8�A!Z����Ds<([fdy��+���^-��S� k�#b/M���cG=�#;�a�[:�Odڣ.XB��X�V[�p�k%��n��.���ڰ�Q��^T�]����h�lF����y�`B���A<��QߩEk���i��2���ր�Ǜv 5��wL��q����%��5Bg���qH�6z�NĽ̽�}�W�����0�Y�)����-���L�,��	]$H92������=��Be1=x�^bN�t���#@Ղ#�^�g�=^I��ӈFm��z�v4?q:�_��O�1<*�es����gPW�,����g4m��C���
�foAE�[(+����0��Q�>���r��y��5��_��!��Õ0Z�#��z�3�㝷�M6eu�����E� �b���+��v��aP�l
O�!�`_��"��;8��6)�ʒ���
�����E|������N�5�Վ�K�~�r�����|L�Lq��<�wb�`Y��E�+-�Nǚ֘��>��>��7�Q�i���n1���=	���.k�z���g�؝+�]�T6|��S��*w��j�}l�8 Y��G�5���U���÷��!�A/�e/��!�I��>��vOU�4g˅��Q�>���O�,������<2��=�^��꣬�) �@g#��kdLݏ���(q{���+�@������[ �z��$��{��*/���� �9��C
Hu�ʱ�cCi]�e���I~�z������c��j騌�����b�&������WT����_�E<OkE�t�)|��	�����o��_.H�.F�_l<��q�z2���vǠ�J�I�7�Μ�i��wXIg�I;]��+�>͟��"=-�-�\$��?�l��v0V�J��L��Y@n��e?�_ �L��e`%.�'�2R�+����]�mc�N���D�C�ۏ7\���Y�jP?�u	��H���s �r��Ł
��nW"�O���B�1��qj�>E��7���-=�o�xU�SO��V��R�r� C��R��T>";n�sL5�=���@���YFř ZD�t��ƥSX�<����y_��B(V�̖]#E���w|�JK��γ�k�L��Gl+��PA��d��p4�'3>un�8�b��V ]�h�q-JPȝ�ܥ��D��A��E���\��	��׮7�j�j��=8R��[0��|�
|��5�R=�^��&�N��%!�R���OF�9m���zִ$��={FD��%L�J�\V�gp{����m�V�.�P�[V�p>�wU���,�V�b!9�L"vPDJ����w��?��Rg�vl�Q�C<�Gr��p �{4��;+S�/!�S�+9U�ĖKW_�pH�w['$������ ��x?:��x���Φ��@���L\İm\Ŕ��t'j@��m�<=
-Q��	��S��:Z/�s�ǆ���9J� ��x�}�Ы�=�N��ռOV!慾݀L\bn�a�OBNo���ė��� e����ܢ���T8:��%.��Hlf嫛<ul=ȭH[+�a��ݘ�UJL�o������d],k�z�Ϻ�9'������,��L��5�x��h�&:����>�������?՚�bE��Jtٺk͝S��"�٦b�J�z*tK(��Ԝ�
�ڎvm�,��hd���vɿ�WH�R����aФq��r��������i�!^�]o��;�
1
6��&KZ3�����щ��)���CU 
�=����<����d���]đ��d1C��E#v3���u%`�PT'OEC�W�<[��vU2=��S)4^w�b���X]~�=������[���f4PG�H�����)�."K ��u��8����W�o� W�80NG���P�0�]�n�
�e�25��J`N��q�#�d��5�_��Y�&�NXq�iӟ
������<�)�}f��	s!����g���{o5�A�=���Ee��C������ĳ����I$��X�![��ݻ�n�+##����Ɍ�%O�:��6#n.Y�i�J~�נT�JH���	t���4&E cL
�Q
�K��AI�&G(Q��Zh	�m���9����a�Μ�jZAu��П��
�#%��=(T��>o�ֿwS�=-z&��~���z(���hp4b��hEħ�����������h:��ѽ��ly�EDH�n�h�[�=v4C�R�/��H��B���ʠ��N���$
�~)χuo(���R�����<��"�	s�ߨ#�9ad"��� �[O7���c�(ř�iP�Bbu1���)fQ�!,���5�A���)�����T��I�)~]���?�ⷔ��y���3`w-�p�}L�����ވuG�C@���S͇�<>o&����=�
��%��fxG�]D�_ @50��vl@:���;2�m��z�/�n�C�%F���\���!�P8��c�`4�iU�-($�܋�� �%ه*) OԺ���#�t�������O1 ���cF�V����3�Cʃ��$�#�FE�(�S(,+����0��p��Ov��|)��8t2`wHh��_�g9�}9Wh�޻�N��=`��6��'��a��k��5{x�-�V{s�݅oVW9�e�^���=��Y��������W���������r_�C
*o��+��S��6z8_����1)�^$]� ��|,M�S�'v]p����ΔD-��y�T;� ��K<E\��k쿖�(2��	��tW^�W/�Y�3D��a��+��e�qUK"�\��fARQ��y�
��r���gIK+k��0�&���1I��G@.XN����10Kſ��^k�݊�jV@��Xʸ���/��++���
�/H��*$`��ۡ�l"��P)0z�#/ٴ�uc�
�}�c��n�)�Ksp0��d�-���ib(8�K���s$6��U���ᖧZ��u�z�K�+����c�K�6W�,���v���E�����2���Ke�-�~�Eqz�N�IaU����A8#��0hT����QJJ�@D�9M,9wv}�9�L*��Z>���i���B,�@,g�cA	����!���¼�q�x�!%�����F.�ˋn�G��pQȜ8>D�r��L����Q�Y��.H�2QӬ!N=Y�u�[�J�@[Ì�?R,n݌�?6��6ET9�>��&ؽ��!���u�����^}�2�����^^ס�`e2�
�����J���%�~��R\�c��[���E�Ƭ%���ѻ�.>2�ݙ��CR���O��Q2V�?��^�rJt����	��M̣�����F��",O���8{�8O"����W(�hp��-����&c-����0F}���x�p;���'VǍ�
��+J��N �}�RIP-
R��/��#Н���eQkgt%��a�j!r{o
?=�#}E2�{^��?˯-��\� �	��?�C��B���s(�������7�0�\�V���n�Ms��LD�D Z!�a�8+S�V8e�D�E�!�EJ�d�Y.$
�+L@�&�(�-?0�p�Dt���&���'��ߤ?h�����9T$�T�F�	����
�����XU'r�[�<���E�L~�'B���J&�K6��D������~�֮��ڇ��t��Ek���Υ�c9w���!�l�qA�ݬ�*�	��ߒ�*���Z�j	0��==�"�m����v�>�蔫��%bǘ���F���k8�����m�:3z$� �7�]���΍4�>�B5�ו���l�F�&2<�oM��P�����Rl��LW�nu���i[�2���Z��� oZ�6xޛ(r�|Q���h��r�%L��\ p�jb�U���%�C������`}̺�-�ʢS�Sd���.�����`��梯�:��B�a�=.�c�ݦ2�x@'���:�4./�E��Ud�qr11ufs�$�/>��p�5�
`�ڒH*ǀ�=�\���+�R24��'P��S�L~�aQ���2�(��h�S�~��%�`��*LiT���B�%s"U�'#���NK�:�h�#�jV�;�._<�&S��:#0ك�g�(��}��Sc)�`R6R��g��hT7���g��3���W��(�|�0��6�G�C}
SvJf;�ڔ��ܔKұֈ]`�gZn�J��)��&�\k���*�F���>ĜMo���y�P[���t�2�F_B��w�v�O��w��*~���Ԓ�ѧ���� ���̍dw�� �a�"�I�<TdD$�8��#��O!���>%$�e�a��!�g��CF��)�̳�u*du@�5����ŝ�(6	V�ZӅ�4�G� �S���Ѡ��G_U�՜y�C�eS ��1	� ��lH8�W+�_ꍦÙf�q� Vć(42�a,��-WGQhE�|RT�����b������u�B�=6b�Ǝ-lqV�-��$��<�(8�;�Kd�H2Jg�o��㎿2�%�p�OT�"�>�;�$������%��gD)��>��c<C���H����r�R����Kv-� �3���@�М"Ġ�1�#�ڐ�e���Ǥ�}�*������3���y�����l� S��b>)�c���]�kɥK�}���4��m�4[+,!�!QϚc�{)-�M�=v��|�Z�F-_��wSp_WQ(�z��d��݇�̙�1M��z�ȆR#�a�6��,��2�בq�>��OW?1����	Iܚ�ӕ�1����K��r#���Qq��.C�YO��~�~��8�4z��Kۚ�G���n�!��l�~a}Ry����4��R+b&{�?Qe�"?=�@g��e$��*�c�RWގٜ�F�*��D	3���mɆђ��J�anf�u�	����5x���t�Tq�p�c���/��Yn��� 3��g�P$z�nJ�D�FJ@R�����uM�G�\��ؿ�K�,���%�j���Ԝ���k^�0V�>����l�v��k�Ƿ����NL������_�G^��d���U�~d@֋vh�+W���緙������9�6c�LfZ��j�~%�/��vua��� 2�\�.�O��R��-�P�E�� �+~}ĺ��R<�g��h�7�a�WV4�Nr%�N"0�~p�6@�{�O�W�?%��=��eSF.�n���`{�1(�W9P$1u|���%V�T���}���z��u��N���U<��P���m��@]�k�����&����!u�r#�ow���\Gw9�Yu$��#|�������F���a�,���c�q�.��?߇^XZ���o<�+��YH7����`�M���	p�6�e�w��kr	�wP[����S��9i� i�"0�;��ݣ¹06�9�tz��&��Dň*��ę�ݫ]t@����x�dt�[*tG9F@٭���r�~CG%��ߋq>��p��gk���C'њ^l:��J����3��V�ר=oU1h��q2��O��_�(�W�X��z�:����EC�R��A�y�D1��N���=�N���ۢ��.eHu������cA�\6�׳�B��
�Ϧ	{G�Ro��+d#i0A���?�V��-	�	δ���hU h}mo�(�l�O_`m9����Kv���^ ?ⰶ��������M�',L�R�lì�|�kn�����tn��v�ө�Q��
@̇6��?e��Я)V�n�vb/m	^��ZL#?2*���u�l릉���WJ�?F�N�d�y�J�Q��E���(d~v��p��W�P��_1�t�e�<��<r݋�s��a�LS(�-�ZV�єKgT$	]�uV�� 4��ƍ �a�,����渟֜�淯ONyl�v+�E����&�|X�>�^D}�"��\�o�(a�фmB�Б��T�/��:��i���ߪ�32���_��{ �+[f����j(�+�������*٭5�oY [fca�S������$��#��Y9jwom�·��}�v�a�f��ULi;[�e�k@�'c!���x>���!�+�^��Nq������*�B;S~=Z�f_�р+s�� ���i����;�ue�f(R��.�%}�aX�-��qB��'���}�~�-�|�?p\ e8̓j�I�~'3Y<t�H,�>v[����ʓ��q�iI�8T��p[���O� 5��Ν�Hv�7�����ɠ���Z�)xIK3�݈��j~i�Si�Q�-�A}�����{o��~utWd��3eWсǚO�*S�)�5����/���6��)��a��"����	������z���� �1�
�ܶ�/��m�\�p|1��Ea.�EM�?��Ta훕�%�v��4[�l&�c�;4fl�?3[֥h�@|�=y#���8�� L2}��R(,��W����_�pS�1[��$��&����߱��(���D�W�0 ��L��9��Kr�Q��(Ee/h0S	�-�Y&�L�vO�08@��M���9��5z^�����a}�mc���;��2$��u��N8�G�������Z�W�be5Q�0�Y(��cM�ejw��}�t¶Ku:��lE��tV1-�� ��T���}����]B�ƗP;"�x,Q}{ט3�.��y(�8��R2�#;�di�B�inG��L-��X��"�'�,h��zG%.K�1��ŌX���*#�2��/p�	Ӗ��o^��ȼ��d�="��AC�����1e����tK�1�� �s��q��D�/O�F �p:&��p���F<��O�8��fWC�ݜ��c���<��C՝H˧�4�J �&\�DX\��V��.!��B�׶��[!8�Ț!Wn��ޥ�Ș��D��o�>g�dz���.G�F.�d���
�������%V�^��8o���;/3d�a��>��BY��ІM&�Vs�N`.��򷞡죴��Α��va�E�0�����*'O8	M�����T����o�j����c{�ڑhf�UNѨ;cΫ�}ޕ�{���
��z��b��BjFJOM�2u�h�{m�.U��k$aG�d��gQ1�Q�|���1����@�3�漣C��Ƨ��P���ZD�:Rn���c-Ӟ��StpWmɶb筗�4�ՓG�ĭ=�34�����Lr�;f��n�Y8WQf�
�&���)K�i
����1���$[TkwUcM���y�o�2����~DE-0�#�8Q�|W��6«�6;6QH���#��&/VC2��t��E�/�h�v:�+��Iҋ2샱��
��'>RL�v�ȻH�q����@�R�X����c��1yD"x ^�S�N�!,���ĝ��8�{�ٜ+��x�|��yCe�w=�<�p���{s�Eù��7����U���x�]L�Vr1��^���n����~�N����\����'2���9�׊���Z��y�=ߐ �EH�OcL��-x�H6�����h��3�]C_"s-F���dٴ�dn����w��&�tj������6o	��E0Ϸ�l�u3�9�y���F��؂�#�2�F��%�(�u>肿�f'�'��cg���ڦ*��
Uj�P~�e��!T��$T�c�,9�ܓ��Zߗ��ՠ�;ehL����.�-��k{3ZCp9�1�lB�4PXiZn�׈�#��a�
V��=�Hfұ�aR�(��QUW�%��lv����s�O.���6Yy$-�:Q��΅߇��/hu��'�MU���B���V�v�므�����#_~:��������*_�/���k(�6�Kf�D����ֆĊP5�U?=��6u�#�<Z0�,�t�D*�и�o��s��8'VA9j�w����i&��{����i�I� Zh+Q���,��Oڪ}�%���$����P��獮���U#m�*I�\��`��W	2}���Kۧ��y	�P���%��""�qk~�U����,픭ct��`��Ƭ���s�k�$��\�y�)hJhCI�te6W�"K��U�(G��ڎd`��.��<g����@w�_�=�u�H���}�in�I�J��VE˶-`�F���xm�:?M8)s����5�Я3G`䝆A�;��Q��J�#�*��?��:c����Y�,ؙ*^��|T�|,]� m.�B#ٯ6ۦ��l�5b��s�����C8� ��]v���A<^���K�z����_���g9I�w�G�m`�I�@n��O 1m6㓎W�1��|��+V��b���K&l��*H*�4g��BDD�I���(��:Pr�M���NDu�B-#6�Դ��ޗAN�J�{�O��'Atdw�H���ȭ||�R鴮c�hIM���ӅiȬ��!��B�[�㜆�#���_?uY2(a{��b��ą��x�8k^PzO1?!��Q�G��Z�*T����,�,�����)�$�2\��8k�3l�A,s�k�� 8��Lq���k"J�V�p�3��3#p�t�-x[鈚;8�(��±$,tw�~���^:L���^�T�+v��G'�؉	!��ٳ�V����Ej:����><�9u����M����z�Kㇰr ��M�{[@�G�+FN����c�@{�# x�R�U�C�M�lچ��+]P�f�\.H�N�a�����L17Wd0�x���Tx��zR��x|�DGSӍ5H+n���!D>�1��s�.�r[o�����(%�)�}g���+�Q9��� \Fb�nN���^U�.M�ߡN��2�:���)�:Fr�<�my�ɾL��J4R����O埆��)�g�����g�O�X�8�Cu�۾E�T�=~�C�Ż��@��_bX�%�S$��Y� "h���=̨j�����~/����l��('(׊$���`�7+g<�{����a��(�f�Ūk�������_b3���~��.]�7��$�G��-��q����!���6��K�u�_:�'�\#p���$ɉ������J��ފcv�
뾙ͤD���aT�cZO��Y��a��\?�P�]�ߡ�=��)d����Ƚ��oyң��#��-!��w��d���N��M+��ĵ��p��z�?.��i�=R�\��Z��:@�7�ْ�����w�������1(��;�1��_��`,!C��zh��	��27�f!��u�J�W\gq�B	�D&�V�Ł��H�i�ރ�T_��f�Ɏ�߱��ml��X�y�¼�/��\4i���}b�Vt�'1Cz~��2T�G�5�'x�_��.�Oj5����G/��^����pc��@j�Fn��o �w!�K�T�#w��/8۳�	�ǘy5�Z͐/4��J�{�5`Jֵ+�d�Q<������h� s��H<�n�3�
+1:��[�
`�An�q���&�-��[�L���̈�wni��`w�G���0�Ԕ7u���j���-QN���\��EC���*���"wJ6ܗ"O�$-~r����aeu�O�/1.�+���y�Q����A�q➭�|�(�s]���h�qU�>V�W�ʔ���r����Ri���ݥ}��g�ս�]g��.����@;����$&M�&r޿�I�h[��KHV.�b���)k��zkEzU�M.$GS��N�ؾs�YD�t�#aT2�G{Q]4U�$�:~��Ǘ�C��_mob.Z���Y�,vbH��A,I���շ�$D�X����LM�� ,9GO�
*�$S�镓9����_<�e�|617o�=I�$�Bߐ�[����l�Ω�g�n��(q�'������	a�gݼ+�~��'����r��K	I�sF�/�oӱ�)��{{�rn�̊�n袍�)V)�GT��^e�V���kJ#h���8�|�Q���tU#5PĢ8�߃d�����58ͱ�֘p�Z�?�ߵ����7,�O�yA����۸-��V,t;�z���ބ�B/���}��+\)��ۼ(�M�NV��6�^YSB�e_?8���5�T�,��-��MWxحY}j�Z�����{��/T�b���u�t��3w�7�Jx/�5��	�����T�+���z����l��41ʺ�X��f؁b�_����LX�����7Pp͕�y�45��*Ixp��@�F�9�	L�>��;�vz��8�8���QaT��#ty��-M�6<���xo��|Xp��8���Y��;�y]3Y���z�T�Y@ݦ"X0W��G9�6�Σ�4�X����"������<Z?t��4s0��d����蠓�,�l�����_
U1WI�ٔ�4�����j�;�h�D�z\ ���T��_��K>QQ�� �R#�t$�},˞�b �%���>s���s����;��ſt�{�|�n�`�<�WH��\�2r����a� Tʍ�z�7(W�5�Շ�sI?&k�}[i�	��]>�!�?�C�*�T�Z�s��v�(1��/K:�B*I!u��cQ!��0� $��-$ޓ*+Au ��;����N�$`0ж���jW�v&�D����{j��F=*���BC�|n ;�(�aE��t4�@���"�z^~�hx�?��Q�*�����dD�/6�"de���U>�g�P)�G.�@Di��F����30c��xm�+�:e�`��4��K���(���Ѡh�(e�%�h~��P���P(#tYڎ{�y)dq��^����	U�r�H�{t�1��x��V����Z*��[�v�43�_Rc@�^��o�oa��w���X�mV3���}�_�������=�A�t5b�o�L@��'��u�^R?�R�&$�82F�(`�&��V:���/�
��љeIiZC�I�	�^���>��E�u��iL��G��<4��Hw�%������j�ȑ��KY.���柔�B4�E��N���&A
�Ղ`����o�)�:�3�^�o�K��b	x���'�����$�x�o,k	[�8<S����;g\�\�w
�a8�� "	�{�(-�^kE���TQ��%n�Nx
5s���s�d�	̰Ȟϯ�����G�\�Y��K��l��r ���c��D��(��kA�@�X�[#Rz�ͫ}j"�����s�M"��(�69Ŗ�o�]٫�j8h�	���붶D�a]���1<R
��!^��bx�w0(����M���̓����������Ű)R{��Bo����=��܉�������[H{ؑ���j��tR�H�M:"�Y�B����<�k���Թ�t�p٥ɛ�b��hl�/u6�+K�x��"�Y7�Զ����v�ȞQ.ҬJ����@�d�-�Zj�y��}��*���~�螪{f8T���q����%9������8A<N4U��u�{��]'lצ5�M�J/di��p���j��4��:��$���m�װ����l����E����k�+
]�������Pl��J"��Ǧ$4�A`X��z�F ��m��|k��Sie�E�����-��a��DO�|b��ll]�
�	0�:\m�I𞾻nտQ����$�_�E@sf�� �w0��s�^��kÆ4ݬ�j;����Ig����*m�e���<���g<_x��i��y;!���%�����z�}hY� J��h`꒞^��ȹ+ڤ`��bN.wnj�[��Lw�ǰ@O&�'cq��w�������/�ַi�]�~�@��I9�t�2S�	����M��>�:im��3��z�r��ͪ�©"��%��,��|P=�:k�g�k؂��f���"ġ^�X�!��E�򾘀��s������u��4̢a�>Q���x�C��~焷�6
�	pTF
�T�n��,�1�
%��8�I���s
ga³T��1V���0��ǀ�2��8�.i<z���D$�F��3]ݟw��8��#��L�J�J�+i�4A[>���|ۨd�U3(�6n��"�ĕ3憐�sR╃K~�W��R}�OY�<�PP@P`���T�$
?��w��|�doU*�p�h��K����hcJx���=�)�R�)�~]9�q���3��oM����11��$!Y�3G�����q5n]������v�<Cm���\��<��k�־Ϟ���FZ9¬٘uN<Zʍ��q�屚�X�����[��)�&�ĉ,@�5l��%��F*��3B���FwXDB���`R��Af�}e#�G��}a��rЦ*z ��j�H?(�`Ş���w���ʲptZ������H����
��?�����[�Ð*��'�k��e��4<Ct��U��H}�@_Y�v�F?��,�:x~�p6������޿p�Wd�����P ,x����c8�蜔���L�g��1W'�~2bp)j��K�_����1�E�N�1�= ��1�z)�����DUo=� D����m�d�/G4\��i��|��7����P�SxW����hDjL�Ffh_�,9;�yN͞u*�`6!.��y9�4�ԡ����'�sqX�2�C��?�#���R�	�ڨ1�����\k�֫���oe<>� e:�\+:%�x���B:�7j�e��OL����֪�{��l�������W؍o�GZ�{�]v���� ɀI=�
X,4IDW�RD��p�^�xWP��SE̼�Ԇ/$Mu},P�H�ED�j���K=�kT{�u�s�u'��#T�0[�e��m�f-��	�[J��r�|�ALcL��획N�i*y�e�v��g	����Q6V(�wU{xB:��*��� ��J�+�������T p)!�<�8W�#F��&��k� ����_pB��_Β���'�u0|l���}dw����B��f����ϫ�K_pZ
WցB�#͝��d싳��J��0ō�J�m1��M�+C��	wǺ��A�,݂zw��c�X�*B�r-��n��%ή�u�*��~nKz��CbNEe�z>@����=xni�4G���F��ME5ٰ���;���`�t<������b6��.�H�Y+AW6s�u�*lc�U�p��O�X[�	�PVv49���s����3J$���\@87�� �:ɢJȫx��L�(�v�໭�AP��ˠ����r��R.,��`�׺��y=�A]]���Tct�9�5$����A�Y���t����r��Pe�u4�#n�/)��/8�c��}�h�����\{)�lYڅ�3"	8�򑅩]*J�:� ��Q��d�f��Cr�؉׏��!�$Уu���*f-��{����ӻ%�Ui���T�	�,�/�r1,��A�e�a�a�� ��D'�9oṣ�׍�Ϫ$f"�Ϳ���J}�h���I3Fk
�}x��J8�
�3�H����^�
r�����x�,q�/ 8�&"����{|ՈFat��M�����0k���]I����(Ԓ[*n�d��l.�t������(��P-����j�� �$+�u��m&��9�l�^�u��؅�,d%b��9ٶ�=}(�G[���eڙ�>G>�A��/D�:���T�O�pOxv�"\q�Va$�'��Сn�����q䰝��b?�C>9��YLZX�7�Dn*���KA[i0H>�]Fa��bNS��(&y+x����{�dCW���X_�ֶu�( ��l���`}gǿ��wa�9���k������K����zI8�����3뱴��Z��8J_($t�wVYFN�Hܿh�������������?PڛwH�R���\?צ0��L���Ƚ�u��t��/���7���U�w��a.��2
2��0�m �qM�B�f�)i%C8�n«R��A�\���F,f�$F�c��K#8X�Nη��p@��F���kk�G~Dck.E�^�Q�ǰ�^	����ˋ�:Q�Ĩf��WM��N��+���36�%��XUl���@�����Ԭ�/�A홾NEB̹���Fc+����.��qkZ�1Z�5~6f1/��� ,9�=��_h�;F��T���!q���PX6�*�Ӥ�є�8�u˹V�	�傿�K[Q�������8ju�B:v0�c�Xp���P��D[k'1�U*q ��\<�v�js �TL��a�h�h�"2!4o���G6���5	��盵�5};{�����^� ��ƿX-yb���L<�@ϵVe\i�4����n��=�|�*��ۭXk^����)������,9��p
2�W�^ɱ�″�X
2+=6+j��b�6�<^��_i0�ye����=�3��dD������ߝ�c/�j���|ȥr��e׼�6���#����Й���������s�%|���T�-/��6�e�W���OU��]�-#�.�e-��Ա繢�Fր�^)d�}�����t�|0���M�Ū����/�O�S���A�Nd?����D���yPVV)Zjq2U|�N8��S�*�~��{��RU�#{�6���ǗLN.�c��;9waY�~�}'��Q9�)
Z��ΐ��������]�ҫ�>�r��yp�0c۾����&�����c</�|e�����-�]�%�t�D�_[�7m���c�;�.�8L�Y�y���eܫ�A%���g���<�R����*-�*l
/�e~ӯ*#mLiU{�.�X�T���y<K�%��h����2���6����;$��}�q*�,�R+�b�:��| ��;�N4	��.��ҙ���Q��g��U�v/i>�8"Ҩu���3q�]�I��A����h�ħ�Pn�@�nK�^�����w��H��;/K�U�D�,���h��������(J�O/�n��;�8�2��,J�nd^+&�HdZb~3|2קӇ�/��쑊N�w��� 7�(��	kH�A�������;<�:�����H�vڈ�8[>�o�,7ڙf��=z"�a��"ȕa���Dz!H-��>)��%�b����s �V)C��P��������Y���
�7��.wtZ�5�6����RI�y���^C�����7\T�DE��A4��g"]|,�?��>H�{�z2kA�r�>�Ȍ���\)T�$��@�.X���s�� �+lf���Y �W~�gqt-1u�j4X��zy��͡�*�6u��?�A�{�Ri4m�f�dwt����Il�A{�@:R�:~5IY�A	�pQ6��shRTy��1p7����3F[���l��O�;����vw���"@�/�9s�S��,*�i�l��OeM��m�� ���W}±�����=�u�w�����_�Z#w ߂�����ڍ{�2xFZ����-}g�S��)h�0�uE��rh��4AM��camF�l��H+&4�vg�`z:�5@,�mf�rޚ���П�l,	�U0+^��3�@��Z8j
i�CR�l]Iq�?�u���My��|`��k�Qe^:�����R|~ {�
��#��t���Xˡ���)*��F�g����غk�w�e*OX�:�8'��?��Vg���
�nj�9	7S�!r�w�����Ĥ�� �*i7�H7��J�O1�J��&�]&�x����F�%��\7�}U�;[l���Q��U+qZ�u�U0&)�}��t>�#6�49�G
o	93_#lSb�&�P��E���p۳QKk�u����@�B�X>���,�$�[�:��%6h׷A	��~�b4�щ���aXvk�$'󴺡?�g�D(�|-C���3tȉ�չ
zmr
'����>̚ipV��AK�lG��z�����hY����D����~��[����&��cVH�x���3ll�E �HcK�m}�:���R����Հ�ʁ�TXʠPaO~������H�uB��Q`��G��n�SG�p���rS��&�B�8��S�ƽ�����s֎�p�_ƈ|���3n�)Sc'`�@$��D�'R}Y
?:�x�?�(K:6۾�=Wݜn�yiӛ� |Op�:����`"c����� ���L +2��������)o�<hqh�Z���A1��50o&t��M:
=�{sO��{ЙXn�E����/����"ƶ{��SV�-D�g�+k�� �qb:g�`�f�PW���|�b�=�P�������z<0�7`SU)�.(�,�r��ǷDL�&��F�ݫ0(<����-�)���pW�G\�k����Z
5�z�'����5����8�q��2:|i�X
a->K;Bխ����Lރ�F�qZ�	�y��8ַ���a�P����7#���Eq�MᶖK���A�Ӿ&� ��m"�8k*Y����4�6&K�j��#΂����oϝ���c����'��Q�;�%����][�CRY�^���O�;f�C��ֲf��?J�I,>��/����>��9�R }ϊǢ�-�bk�$1q�ڍ�c�ѵ"��b�o�#Q6^�ֽ�]d�\�`j��6�4��1�]���V"��M� 3�&�$wJ�G_Ψ�JS�HW۳-�$~K�`*�����s&���Qsj�Y'?��g����Q��!dڍzq��hWВ�NbJM~���`\�n��.�Z�z��Ƒ3V$}$���/�RZ���p�Y��{��vm�}9h�9�
�υ�<����3�*v�̳��V(yt_��)P���Pq����XuhR�J
H���љ�1�p�"�^��l��o��>��%���`eT��e��uʹݎD��"������ڏא&�M��hs��h��>��tB�H3=(^0x�N�u�����嗺�zl�ئ �;;N�U�b�R��z�T��'�j��cb��!�@ܳ0:Ta@��oj ��!�w`������bq`�����7��5`+�Sh�re�{���é�ye_�t�c>�ֱ3|{Vۅ6�e�l\?i��Q�����[A��#�ħZ�HDI�9�U�gf��3u9�<)� �:hy�=�vӤ�������n�[G_��`	� 4�D��xX���� 7�JvG"=u����M�r�f��&��|xZ��R�^����F��ݻ�c\�P7�wM3��.�R@��=��Dj��s6/oN�?,kW�.k���޻���n�^��6��D4�U��Bהɧ�~я/a1´�����W�D�x�����Y����`�+2`ȩ��YN�0���_�
�.�8��<����2�`���hI�.0T��TO&�'����Z3dxxՋ?	v2���C\+������̑��p�������I!���]���EJwMW#�V��6���;#`Tvb��|M���+D��E(y�m}�$���5Zp\��i��=��+%�E6�氿�{��,,�#~⦕��XdQ>�~�����8�:����y5�r<s�s��nj^I�cj�����O�&�C0A��o�s�bm�!*�+{<�Y�р��6;-�4D]"僊@)�#�u�:�"��7��k���g�'��}�_+����)/Ό��ت�󛱪��S�O`�N�f�͘��G�Nk��'|�Z�<hR���]�~�SL�\U L<�oPf���b2p���f�~7����)�<��é36�4Y�RCq�|Z�A�q޶7�b����38��ƿr^��/K荣�UV�:�f���J5)� /��)�a>��=:,unߗ#Xu��maő<���/����cl��,�Ma]N��!͉�� 
�8��J���/��y��cx8�'�cl�d�x%+y�I�I�L���=;r�*�� .߉���vp����*�����Fӝ,'E�V�n�_�t5fٸ���o�y�_y�y&�I�=�~9�2��s�Oд ���<um.�4��؆�6r��rŖ�ѩ��1
��9c��p0.���qOQ!�c��(�iY�M�N�/��HZ���˻��w�$?�ߠ.P�8�k���%?��7ӿ�B�:x��ơ_N��nش�C�(&�$�IkP	�r��1��R`g�}��DɆ��+�Z"�v^>x�ԇ0�N`�VO�p��Z[��{��|$拪+&,=W��=Z�Fu�,�Z����;xm3��a���B���*{�V�)"��&��e�+����F�yw�<eR�M���Q��*W����.
0��B�p_�G>r �n��H~��j}q�J�� �����n��d#��f�Q��#t=�_%Ў��̝��{�����U�^o{7���� ����Ҋ��^w` ,�����|a�N�T����X35�t�ls#Y<,�M��$?��[coR��v�UA`�,�[N�YB��" {��D�~�R�0<��m�uF�_cJ7l���-UM>VC�hpm�U�����hF|�i��h�e
�_د�����Za��\�!�S)�V�.o��(�/2���B_楐�BqD�}vmVLu����7%g���_)ܿ$�6���%�؛K*}�����8E>xB����ǎ겈����]�b���B�*&o��4�f���+�4���"G��I��V��u(%�oO�.itM[�x��c<����2o��D���5왶.�&�����I�T���6��Ѝ!c��Q� �S�՚k��x:b�aB�����)�he��YZd�H�p�>���|T/?-��z�V{8�6UN
I��H���<
 �i4N��������-.�]���P��p9D��w���s�ك�����(a��sG�'K �ާ[�c�(XM�`��0@�\�����Ⱦ��ɑ�Mr�����?M�\[�1��z�M��d�~� +�y��:�&.x)��`���p��Ffv��Ӌ�A�e�dлb��4�L��y�ؐ텪�iD����_��O��+����a�^ ��w��4N�g�3ْ��;q?��m�G�J�m�F��.���#�t�8�����^Sm���3�����13�@��Qw�ō��7p-����=`� �م{����v����� ���zb�3��@���̣H"¢�M��d;`5�=�l��^}&�J�W�P�\��AF</��ݥ~y��#sW��S���:J�F:�gw�<ʅM�Bi��5����j�?�n�H4�<�\��	1 ߁n��%_��*�ٴ@���Us�榽y��ۤ��A���fZD!�t8��U�Dǀ��>*Y�鶳�};�����[��t���Ov�&�.s���O̿�	8�I�]�q#�~�h&1�8���V�?%�3f=�C?�˹����#6_l�itDCT9c���p�+�b���;��A�5�_ҕX�+��"Kq:�`|��P4K�Qj�zn��=��Ǧ��B�:"<8P��@y��2��g��S����j�<ڂ@=h�|��rq���@�u+i�e�H�_Qf��y*�L�0����s�c�Ω�Ay��h(P��Ž��'�ZQ��v�n�o�8�Ώ]胞nɟ��dO�Q�]��#N62YTK@M����0��ݟy<�-���]l�E�$�W>R�(-�_c��J�%�����B\iѷ��AHy$⤳nr��fa�ĳ"Y�!2b��ٗ}�������;��Lq���լ�bD�EV��0�p,g�?O���d��lZ��ΩU�H�$/�sIt�°�����,����w���"z� HdL-0ђjY�FV�mn�����|�m=�n�sN�	���p��ي���δ����m�8���q�XSA���Kj`0-�j̐;K�	�����'��?|��K�a|�X�L��#+R�mjQH��X�����<�����W�fO(#�r��a`R��
����I�������xB]��[���VI&�l�M+I�"�y��G}�I2&�!�x(t�qP��t���� ��϶��6UHw4�9��,Hd����8WAsT(��E�2�|ޡ��ͮs�݁�" ���qC$j����w@vswU��֞�&�;t��~�/"�ѷ)z<�Qh��g�n���5��m$��.���M�/�F7{���q$9�Q�AC���&w��u\;*޸nZae���Ob��+T��L���㸏U�)u�Ďi��7��e�o����[1���tu�p�WG���ݳ�Y�z�	�6eˍ��l�FW�}�b�(W:|��� ��77v�ZgL��ȶb�F|���3���&M�O�l�EH��k������\|h��k�ϵ�������9���v��$���s]�@�w;�`X�yˤm`��<���?�ț��x�$Ĉ��� ֒Tۊ$ ���2�E���m}���բ�-�0j�4��+D��=����đ;�iH�Sĩ�X�!����q����Lx�q���'K\K��2���,˂�� cͳ��%:���a��LF�*�3Ӟl����vS����9@ϗ�O|��0��H;�LܻQ�ܯ
���6�#3	�̆@s2���wmbDb2{�쯺E��ޙ�b��6D��0�3��,5�Z1[�.���Ir1h�/��b�`���� #LCDƗ�T�玒�oiԛ�B����C#���R��8�r��N#p����Ki��|3�Uu��{"�q��O5<vf|��1�����5Sg�W���A1��V'[*?��
ɣH�o�s�#;J�1c�7�/Wh�$�S����Y9�E�J��4cϋ�D'] ܪ���EU�|�f��vL,gl�`�߼���Uر�����湕ǻ���t��P�dy�9h�zJ<���P`����`�q`}��l��!����?܆���N�.�54Ǟ�s�/�����}�.��mE���6Lw8JE�0�CK�Y�3 2o�	Վm�-g�H�W�d��(a��bVS]Ra�$%�+�Q4qQ#��_嵰̗*�r�H��M��;�P�-�<l�0�ɋ`J��()�]���F�����k0�H!��j��X/�_�i�������,��Hx���_^1��S8��XR/KOf�h��&:�&�Xcg�{�iE����#&M��7��k&[ؤ"c5�gI��a��ͤ��[�y!�	�m[���c��i��S�Q���"`ȈL��M�rr3�g��'A���aMgv�g^�""����]ͥj�?� q���?�i�s&���#�GHPW�d���}�́����A���`(<K�T-�lw�1���K�����'<�zc��Ӷ�5i�M��t����w+�ܳ���(.=j\��*8"ު���6/N�Ƽ1�%f���z�M`�Wy�#�̷L��(�o�{���JP��k;�]ι_F�~9!�-S�V��c.�˭�j�p� ����ӃO�7g3��Cb9�vK#:���~�b� ��Z�U��da�
Z��V��ʇ�@ť�����z$KR����K��
����-�;ͫ�e��g`�~ɞ(�j�Ra��r9Z��:7�����8�|u(;���9�F�f�j#˛�2_#	9���=�Q͋�����Ł)?����	㒽lL��ƈ0E�
`�3E�Q�M�����6y�Zh�B���h�.5�r.��f�؅�/�����*�R���t����dgd+��5�M�ȵ���3Փ��p;�1���&���K��P�kX�5aj1JCP��0�K���%�#&�����GX-=�Ѡ�?d��L��"���N��¹��Vk�S����q��"������]?=���-`g���jJY���QMhkX��jj��u��Pn6�탿��Z�]*�� ��.��\���2�]f��K)��i)�>�E�ڪ��V�3����k�-o�����9�ʾPT:�j$r�.;�It����9�\D�y�*��yv6`+���|pIz���C? �����)��
r���,�Jv���v����D�u�tc��b����=$�����*�o��Y��{�:�(��{-�J�%�oP��}�綡lC��������^O��O�uuIw��6�}�[J!���X�r|��4^4d��M���z�sL�L<�ˤ7EV�XƊX:!�Ʉ22��LsQ��;I��)}g&c$��H�8�Ӻ,0�7P2�"q	,jl|72�P��O⤦�	sI@��~�?`u�o荋ȱ�1�n����/���F�B��l��ݦj

_?5E0��i�G�|Kg��=J���*S�n�I��b��#t���*�R
�\��&t�N�k���(�HYdb���𑺷xȖ�κ��W�e9A���
�ޛK�z�wjz����u^�fR;R�`�w�#Xzfp�\M�ԚGdЫ�������X�r7�����
lKăAK{ݴ�M��GLBW':𡣚�ᑖt?E�P�x'w#9L4t�P�џmE��+}�?���0%PI���6T~t����;R�5�f���{�FJ���Z#�iz��0������Չ�%*�\�I�W�5�&��:1c��pWeb΀��𼇰�Ƚ���ܗJʼ��g��m�W)l� aQa)��v�)	�\���ĺ6bK4���>ן(�L{[����\�"���F�bH���%nTh���n���4Z
W�~����G�V�֣#�3��u�����(�@E	�w�6�0Y���.G�R��������iyc������I}L�NÈ|����@�'p6Ӎ��Z��b�S(��r=�;��'�ϿM�X�̦[%���N/��1�]�eRT���s�(��v�04:y��|�~ο�lbek��P#n%�$��ݍ�ӻ>���a��3Ì-hesUZT�� �`����_(~�=��Z������.,D����1�il�V6��@�[������Ouysɹ��ڟ�~�7Rr}�4�����䡜��+���B�5m��q�h�ҿ7[n�]�ݯ���3���s�l4��3�!g��p�5�\e,��k6Xk�n,
���� >�� �x��7pU�gN��"��gAAV첔֋_���n��_H�`�!h�Z�N&J�i�����C�P��h���c��S�`jM:N��/�7O-)PW�T���LsZ�Y箚-4e$߫�#�hw�Ƨ�MJ9�(�����qaY9�M�����Vd��{�o�AQqZ_�d�-F�D+������P�����0�{Pjy�ֵx�t�RD�ǎ[nϷ҆ϢKK�a0�N[w=���s�-����EHe��/�%z9��ٙ9�V�kob1�S�i�"���K	���K�{�}��j�2S1������F5O�'�u���;�o�O_��r�EϧV���&=ꡓѽg�2c�$�G�����*g�H���,1�ˠG��b�[�Ge)��8�P�h�����b�\����6*׺u׏��aV�'�Ĥ%�CZ`$�ߓ{��}A���sk�#��m�ObT��Z�cd�% ���<�4v��C:2�[p{w�T��L��#���{*�4�)�N���ç32u�<S��*�l����1�Q'Km5� �OvL�cӷе�j}<����3�'�%��uǿ�:�O��R���÷��̛��$��P[`����oQRR����6�����Y���6�������9�
��j.�ND�_��������Q���G�Psjb(g��5�3�3��Le_K�����^�V%�r3*G�3�8,30���(�d��2-k��l��B�_~/w������LB~t�3����T���"&,�����>���C��LW�[��{Ti�m���$0T�9��h=�܏�6l�L�Z��C�����QM�"W^��c{�|2B=4����-��!!��1)�s?�����wC�/d����w���l<�#q.�t�8
Uf��h'gj��FK�Q�ne'p�1w�k ؕ)�(0����#���Er�-sW�ջ�}0�s�-M��m�����yNQ�������X�Ó)K
�]YwB6x@Z�?�����'i�ڀL�C�v�Pi;�����	7oo�:<	��m��J�/q���U��z���{��V �����8N���J��0;�\���6��.v2�D��4Q����>AH�1��v�*">�Q�V�}�y|&�/�|<Z��+�l9�Vd؄�A��O]�rI
�����(_���(en}�<��;�Pb�SKmR*�6�p0��0�/�"V?�{�Ș��f� d~@�[h���2\�U�qk������y�.q�h����O��a�X�Bu��Oh��:�Q��l�ᏱG���k��g������ ĕp)�4B����r2oN���&�Qjc��a��}Y���w���5���#�|ؑ���!|��sǱ��u�b����ʡ��3#��/E�uu� ��tj&=l3V��~��0A�o�P��E�h�8��dy���-�R�Ž��Bu�� �;�)���<���U�G��A����L��g�C8�6��A�J�ɧq����XJS�X��Jر6���0��.u��W�V���P<�����P=1�_2w	Ż�jE�a��#�?\������@�DtJ�o�ǹ����<<�;U�����O�|�MyX�l�]���P	���/��=B��օtQ��.pF�:{X�����Bwf��dF��#JÌ7HP���ih�Q�b�lKH<�Ҡ&��8z���sB}���d-��}�4������A��F�G/d/�W�WO�pR����Yч��������q%��	�G���X��ֹ���z�>7�%�-N�m��`?L5���w���R��^`R��*�TS�"Ȟ�=	 i���K,�C��N�J�Wۓ���������e&A`~�~e����F&MR}���/F�m���a��Ua�����Až�z�{��1��*�G���C��8��������XdO�mЙ�ř�ˆ^����@�<[+m_��	0y|�o�҂���&c;*��~"QX�
B��%��B1Yo����PS1�wBB� &L\��a�1��`����4��uA��'�c=?:�Ď�=#tK�$�^d��ː�.EBl��Nx��v���G�Ȁ��	u�Q�Ày#����_8L���9� \�ϛ$/FW�C�G���K81��J�� ��osNa%zWn�"{]���|�%ة��<��:��]Z�ݤ�.}I
N�8���^������ui�ʞcw�z#���S��h�J�("i��I����l�'SOv����.L�N�GoZF�mP$�guF%�$�=t�ܖ������s���
�H�{RI��k^�� .O&-`�\�/)@@\�Zl��8k^Y�����H��\���4����M����s_㲚�t*Δ��\�X ���5�L��؃яO,�f�.-��b+�-�F�d�
9�9��ߵ�c�n�|��*���l�-K���w@>#ў���n�'-C}�ǝ,Br/+g��t�3V&6TAP0�c����l?"檊���Njǣ;��W(��'�|Q�k�Lbu�w�霑�c��cB��� 6�>T2~��
��zQB)�9J�٢]j���_l�-�%ʀ���[�jK���uL�*,�`C������'R�f.�*'�{��*U��8ĳs��f<{(�$ {f��z��mT뢄��� ���4e(}�"�wx]�C-��gt�-� �ΰ?�<���W�`ƴ1�� c���-5A@�����bWx�g����E@�e͐�ҹM����������e���i0�p���UJ'���W�2Z��)�r��ne%�h�5��6�5q}�	���Ϳ����P5[A6���ȗ�|�h'�u(nij�̳Ue��]S�F�¾&��tힼ�t篝Pv�WV�i��{_|�)Œ���E���.����e���K�@�����r��/? ̕��e��i���
�(�$�\��炟��[��Y���Y��@Ȅۮ>Ќ�P/��l���N��=�+o\�{r\�{���Y����d�)��]��,*���q�W�Ko�X =�.�I\]��;�� ��mX���ɑ�nWE�?����93�]q�
��X�^uN�%�M��9)�s/�-���P�'�"���`M�0��4��G"Y�Ւ5�`o�(]g���:�x4(�ؗ$�`M�ӱ��T���eg�,!��l�-�W��E�tK��pR#��G�.{�j�`,TA{�sV�����mŅ�X�^�nD��j֖?^ÿSUCJ៕�8��5c�����/�i�C����_�'����@Na"�w*�_e��h#S�];�x��f��
9�*����c��c�b���.[���zra���VN�#�	&����3�K�:�7��_�sG�@�����1�h��q�	�*�
�����M)�Z��������B�Y�R��1]�5؊rfq��e_n�5���=ڭC7[����RL�*������|l6=�㡜C��_{
�b"Ng�_咱TY�=���0/�?��;o]��	�f�M
��I�����[?�@x�5�!�y��O&�װFĕ����9j��^W�Ǖ#ݣ��خ����Ӯq}����ٝ�ƍ����C�)�@"�/yC^x���M���翶��kC���:u��3��"\ĩ�����9|�d���q-��ٺ��Qۣu%P�=�J�^zk�\�Q�Q��ф�i>"r�:�@zi-�SV��@�-�T�Nw�|��O"H���=g�bU�2��Xx#�� DNv�Ps'}��<V]�e.W���&6deڏ���
M tk~mM���x�.��ȑ�GX�b��~���B����ܶF�]��� @z�� ��1�pɞY��a^�섞���π��F��7-�Qc�y����@t0���J�5�.����2�6"��� ��"W�#�#_��ē����	��	��G~}��!��n��A��5p�"�D�D/؆��Y�Ό��u�k���z%��Vi�Wx�|����5u����Ǒ�s���L�h1����4*mRGh�2�"ѕ_iaTY�~�N�{�k�C��!#ۈ	7���}����=�M���e�&��,w�\	�/�aΉ�?��T6����A�p���w\��\�;eq��\[!���]���-A��+:8�E�?S�va�)';)����]羔���E���r@h�lW=�f�f�k��Z����������1�eYyA���IV%c�$$�S+x6;�����}h)��;�+(� �V5TL�)�{���ʝ��9�ު��92�d̸�Y�i�s�Q�<���7$՝wv�t�9=I*S�W	���t���b���xh��8a5J�����)�~%��[�6d2/��bݰL�eW��ɭ��>��P6t�)1���Uz��O[�'��u
l	��Lg �}�/�(k�pD+l�5TB�1�i7~Mtv���k� ������w�74-�F������ 1�bk/1Q�u�g��I�oŻR�.RL9�Uwg�HO�0{�8���6*���:Z�	����z�s����O��!,؞�z�/O�i
n��-G&a����n�&�SU�����Gz�A��<�\?�p��&8 K��sO��9O����Sl4-�[��镈�\iJPO�@R�z=ؔL���闉�D�1�v�!�[� !5��a~�AS
bn|��k�J�}�ܸq�8ߪ���� �;���)�_��N�xl|N3���-�Ö!���CഇP�#�[w#C^�Q!B����� ��>��nؘ�3�J��N�7�%���|�4�.2���3
g�	�S<�'��@��m���t(�hm���@��]���tY�'�~���=�b8��{ÕA*�t����K����4�Rto��V�\�J�$s.�|�)�j)����M�@��� ���F���A�t��Hj.��I�W�*QN�#��
����G��.XY��2sWHio��
���G����|�O�_Dd��q����N+��W�ռy��	��~-�9)w�+꟝=�/���mCm^�m�UG�j�{+��'�2�������Gˇ����j�sΖg����f�	��s����TܯbH���f���YL���'.�:+�r�h��o* 7q���Yo#�-��[�^�c馜у.C,}R{�1�fH}�����D�GŷMiD�5[�ѝ�^�c	��c��z�!`y~�)�����1n4LOA2��}R9��c�� o��R���ڇB���C��.Ԫy�'����{��}E�c'�O�`mPZ����(=�:8���x���߬�a3��b�B}��\`$���qe�7QP�@�ݪ���zC���"�	:�͡Z焭�5���2/��8�J���G��jk�	���`��1��[���Y�z�U	�Z�5����
l�g|�l�	TY=,E�\}�Dt��,�v:}䱬��֨��6<g�B1s�W�����ܐ�6��țT(��`1+J��~jADoE�rI[�3�=�����Mt
�a��χ>tY@k ǰsLog���u�����%�x�`���z%噹�!!SY{�:)笗5ޣ����NI�����{�d�\C,�}:������RJ��wA"�z��
�����A>Q=��VˮMmkgn}m�@&�7m������N@'�'R'��J�o�=�i`��oXl�<��[@�W������<�~��_/�l�]���H�еC_;��,2���3�.�H��*�,�\?�+*Cmɍ�Y)�����η�;����5�R&#Y��f[�h4����[H^��gx��HZk�a�=���YUB)C�-��lfAڛ>q���o㚼a�[����n�TE�&�u�b� �>Y��^ҋ:y��, '��ᳩ�G���8=���Zs&����F�A���	L�H���=��b���@=����r�ʾ<����2I�%����g�[4�U�DK����s��.�[�� �;�̷���x���\+�6O��.��m��vN��n��6�9����!�~J-��y�x���)��	6�r5�vL��*�Dr��O,��y�/%�8��~i����pu�y2�絘`�F�ka�������dc���`Y}�9������h��9K�V�3�I)'��-<��" ��*�D�>K%Gs��E5�
#y��9�Rs��P��?�΁��� �Zhp��c[\|�<PI�,��6��@���
�_���D�^���E����}au��
aJר�A<�rk7�bPmnL�]��ղ��S���U��IL�^�`޷���?^3�v����ir9D��<)[ߣt��}��!�]��SM�(�3?_���l�v��9��u��av�*J<�W��OΉ�G?!|��k	gX`��a�e��(B�Y~���ޮbɚ�"�	��Z���4tX%Z<����R��PAI�D:�-�-�%�x��j|���hVL�1�b#�W`���5|q�(qӆ�BM���	\C�TVU2ϟn�~j\z�7��B��b3���;��X�p�9�\��'�lւ
��:[?�s /�����v��!:l������=�^�Z�hL�kVA���Z��aݜ?������PkT����Gݶf�6���~�-F���P�W�E�!R�ׄ�7��Ŭ;�S��uG���?/(����l���rʱ"ys��K�'r�VM�M�t�8��/܈v5{ۈQ� ���z�K��=��>E]i��/W��gsEs�'��/h�;C�^�Ԝ��_�A%C�C��D�"L����EE���5�0�'�o�e��4��"M���O�>��-{�dX�B�e�Ҷ�A����EQ"�EJ֠k0�b_�/|S�1��6�{�hc��Ĉ�U�az�!��ڳ�(�d� ��8:�nU!�tTH�k�z��͝�6���phv�j�*)ב�8��Ls{.�Q��6�-�,!��c��r�*Qb��1��S��QIH�Ch\�(~5'��M�y%���6
ZH8ұ�)dx!���>Ǽd���?����p*��2�*�H����NU7�
�E*� Փ���0��N���E̪�A�+$�8�J�7]�����k~�{D���� �����{d��E��5��	���1\ ɒ��q��?�!�@a�p-��;���_(t�����d�G�B�(��W�|�U�����yO[v=�
*�������e.&�4��������LQ���>KZ��VIH��N4z`x��Z��맒�+i�WZg�R��Io�Qfk��!;k�&?x��?L�Lņ��JH���ލ�ku�Ѿ�ޔ9t�3xiT� �#1V*�z������tɒ�!�3�1�?�5�k��L�j�	sT`E�38������#���«�=�.�@���ȇ�
�64�sn!Q]j:[?I�O߼�Y�.o��"u�M�eyGT,��v���˚�I.�2ב������+�cK|����UM=�������u���vE���8��(�:�/����n֔��.cFh�t:����(Vy��-0:N��{J-����] EnNM�B�����@��,糾�E�_3L\�e��a�m�)���)�ዉY���;ד�������UoU0��r\h6wx@��c��p�^��H�!���5W�>�.��׺)⪚U����ƕUV�|�U�j����A��R���G;��-�s�%�d���l,�Dwn�h����gv��?� �f6��A_������E���?/(�!��F4�G����X^�Ɗ�G=�Ko�JRm j7o��mp�t*�	f�q`?̪���ًv��8�[��a)*ҊG�t�f0C��������ܱ�6�[��2 T�P����e�R�O�m����WL��=���E��"�����@�D,o`��t}ƟJ�RP��'ًHc�g��C���ч�m��h_җ,=���^�ڌ2Q�)+�Kbi��M[���
��Zabt�g�:g �gEu2����E؀1�&;��CI6@���y� gܶ�?Do�S�6};~���YC�r�g^RP6H��o�j�����z��)5�h[���G���sc>ѧ�B�5s	)�w�k���R���mw��$��&������D��k�dY�O��Z���h@��K`�eu�����帟^μc�c�1#�"��k���y���c�$�BD=�ū�cm+>$�a�U�;�E����($����µ�W�}*��{q��wйj l�϶jB꒖
�Ջ�~���D1G�I{-S��RMn�e����=�ނ&�8l�'B&�H8��O�̬��qzjD~Zw)�Ŝ���Eu̕�oK:Kws�{R����~qQR�c$5��"��%N2�� �@X3 �X0��(��d�mZ�t�4Aq�.c����`Ta������/��-���wڠ���٤�t� *����^L�E�'��������\nw�l/#�<�ї�k9���D��!�Ë������Mw`_�)��`����-�������g�yh�~�,o�e3?e�������0�T����;�AZE!�h��Č�V�t�L�^�a����25~#��ϭW�p=�����Y��(�J��Z�ܴ�M�2������z�MT���0�f����\��O����R �h\V�Is��~���O�O� 2@UJk�H���w���@��>I+n�i��(gW^��ɂ�G��V�!��Q�<�rD�0���v�o���7��>��s�'�n1�3��҈�j�DOA>%{�|u�J���IPfj�L�s���>=�+nղ�-j�I��R$}�H���w>�=�(�>c����@U#x�q���C"�� ԖZKQm����`=΀ �9$K�55҄�qi6�Y�����SB{E:n��o�,����B�GV$�_/+=��rk����Z֟H�E;p�OL���±^hN(2���z#�B�O�K�zῊ��ۦv�YBX�@I��l�v7Y��/(�Xu���ς]*`���J~u�����j����G)�������o�ї��^���*Y`$�&w�����kre����w�1z<�-eJi3֊^Nr�eS�\��b__� ^�z2Y�6�]I�ۦ�ԝ��"��lë����3�c9�pv�7S}��k>�*�$`����V�h&|M���%��e�Z�g��ڡ@II�P���><ܚ���@_L+�� Fa����r���B�:`s�U������ U���6�1͉�'��8��x�h�h���Rr��aAY>-����,�+Gw�G�{�J/�.��e��#�����"$��|�M�4�7f�P<<�����hp���v��:��.cx�{�.��k%��r
�:|����[&�o��P;��x��D�p lD�����mj�#I�t� �RB$����m�P�gk���%�2-`����v�'��b�RQ6P�.)GJ�e�3��1r�u&�%ĕ���eٹ�T�9�c�ԇ�����,��������e�׸y7n���
Q6���?���J�X�4yO��"�ZeWb7�e0�N��T�Q��$n~n6|y��2���`[�[����|�	�ߪ0(�.dc�)0��J�V�)��;50��І��\��5�yVЛ�n��P<#ɍ� 1�d|R�A�|Ą��,�U����Áv��� r7'�ŚzP����&�Ԓ]k��&�l���� p���U|���b
Rɚ����Ǎ�����#͡Lz%u
'�\�Ƈ��W�c�\��*��W�R�ўEd&�@	ҳ&��"�ݛtq�%<ETژ`Z$�!k^}�@��~���a�E�4�iD;��=g~�������Q�$�"8U����u��u>���߄��`c�4�mܜ9oa�-7T^�ǅ3b~r�+I��?��޶ְ;�^$0~��A#��L�j�}���L���(�ľ�h��/096�`:�xٹ���H� ���P�Qf����z�y����փ�g>J9=�aB������i�e?���G��$NA
�	��6��ZNBQb�a0m.�6א}/kߚ���\z�V���F� �<�#��M�*=�C ���+���?�s�f�zd[��w�Nxe�S.ޭ�Ȱ:H��9w�9�X2��k��4� vYfn�����
�L���p���ـ�@z Q���S��� H^h��)�5�ܚ�Vki���7
�e�� ��0���Co��4��Pv���@��鷜O�t�D�r�"�&�x=�j�z���&��Yb5;�Q���>���Vϣ)����~���N�ɚ��Ȋcpe/h�ўel~�ڛ�D�6�V��L$��}�Pb��K�W0���-a����ڻ>��Y�O��|9-�H�s�Yw�(4��թ�h�//zG9�z�#�ļ�*��/ʧ��G������!-���+��S�/�
6t���7��{sU�t��%�����8�dN� &Nm`ZR݂;�M]��e	-�k;�(�n�JD/T�씺�8TL N�`x/��2�'��0��+���cb	���5I6�t�F�P��(�LU�ru 騮���;��i�cL-�Bpc4)ݢ�����6|!��9���_�4��@�s��f�A�E����ՠ.n7�.e�עئ���z�;k�l��7}�>ziA�̥��*∍X��<.���-��j�jf�ZR�@j���H��o��n�`"oc-ٕ%$��c�#L<�[+�v����EL�aZZJ��v����7��!��뾓B�W�U+�)���M��\���� {GEܞZVi0���`�����^�E��5��&��'(��ɱN.�V�'R*� ��5$֐�R}b\[�c�|SB�쬫�Y��o��Wۛ@��?�M�plt�r�����]���αq�+���%�E���S6�*��Q�B�j3a�"�{�+�g��'��c:�ӣ�0�;ͅ�Fm3Kp1���
in<X���'���L��ܾ��};P%'vjA�l�G9Ѯ4�92��u��0y�\�ҫ|,�9�>��MJ��l��%�Y�`�-�z �A%��M%�oo:[b�r-�%}m���dlt3��GY&B����Sr�����y<ǜf�(����K��d��W�3�!P�7Bv$��D���7B��,DC�0�4�C=�N<�S�=u���� �ɔoDbeg��vaȮ�X'��+��_��2����a��Qj���[��1���{?s%k�T�9�,��%�2��� ���&^~=)e��4��m�ہ��h�ڍ~���ni���8�F4e�_�q��.��掤�Ii��#Gږ�X(�Sh�����&��M1�95�AѧmS�H�ɫ��[��E����z=��;�C9����ab�i<2ތ<6���#��7!Qd�ަ�);�$���d��g���Ȳ�ſq�
ٴG7k"A�#hs�������#泔�)���
E�`s�f��)�׆�^���?�\U	G�\/jP3��T'o_#�L�6�a�hC%5AA.@S����_��9�
�������s{�o;���ʹ��)^�ka[s~�Q3N�B�u!d��{f)�J-��Y��4F)2C}��:����A�=Y�/O�{��l�	�H��n9������*��.���Qk:U�guu�'���{�{��h�)n������v�ǌt���N��5�51�W��X�	���A��+�������*,�
t���.�%�]�����D(?���ƀX�8��қ=�5�")�����X����hA�uR�ڊ���|�c� X��:b��`���$��^��3��bz�.�h�o����\�IX�o��b�_L�l'6���eJ\���Cɲ�;�-��<��.~p��ʈ>ΤBJ̻G5��/�Yy�L3��X��q*d�_vZ�d�
bm�]�)�C��Ic)��*/�3P�qQi8��@_�c,�oZ1�1)�%�Sw��ԘW0��v�p�G���!ì��sl>��਋~�P_�HYh��»]�8�
��
��9r���Y3g���}��G���F �w��� �R�G�IfS�]�r^y�}F�&!�Tu�f�qD�*л��V�C�!�B��II�%�����4^��cX�����	�%%K�Z�t�s_ӵ%/��rH���]�{�+�8b��
V����-���շ_����0����
}�JOP{���R3�>�kq^:5�!����l.�\.7�3�4���ZUI1j�.�&vS�.)�=�Z�êܦ�]���ն�W^����0s����Ԣۢ9q'�R���C����� mA�B9<���2�̂��xx����J:v�����-{�Q2��� ��:Ek����g��D��fVI;�v_�6{W����M� ��'u��Ќ� 8T�a��!�%:�w1wI+*�Э/Q)��q�W#��*"K���B���H5�~�T�p����y�����$����~��lH{�B����s�]�Dc�u��}�`�ey������)q�i^_����/�{ ��~驥�s�j&
_O�Ă�| �	�d��Tw$����-��2�뉄7
������Gn������S�M�[��2؞W��B��p����.[��i�p��.s�Yg��P�2үc�/ߙ�h�����5� o�(��N��R���[j�Z�~��󒳍������Hl�`c�8dƜ�P�՟J3&�޾�)f���e	@K:�3�K��Z��b�T�c�ޛB��C�R@�M��'����-��mx����/�+�:�2ǅ �9R��G�Ķ�}c����tl˳���k���d�M��8���P-����ņ�W�X|�\��7��H��V�+3k�u(;+>��I��,d���/��[��9 �AH]h<�kVt	�ϲq.넣?٨1��@y3kzI.����L%u`���:��#��lf.
-
D��ʞFkQ@8P��3�/k�Ò$���T*�S�LO�W�ċ����9�EWC\�w�*�t[��@�Z�M���v�R$Gs�k�V���873�7�5Һ�%,��1bi��X�E�7"�� fLU���rS��ƪ�8[��E_T��XfE������(��C��+���dΐ��?�|n3�;������!-���@9�����_�P~Ɵy�j��i��Hr�G�x���_���ɧfpl���]mS��Eo���t ��S�f7?�b��?$Hg�(��g���c�G��o�)}ze�͖Ҵ�3y ����S_�������v��M�3�f
�H<�ځ�u>�P���X*��߁�g��3�#����.��Q�O�_6_m�7�h:��ec�YY�{���`!��!�G��Ce��[�P<����R�4,@�5�T/PC~+ _JCL^�^�7$o%�n�i+'�/���uW�|?���6���ˏ�����j�.�`?�ƥ��Ĥ�9�����������t��H�O��� �&c���?�
��[(�66`@���_\Ryje�Xѿ�}:r@�aO���h(�&�X3u�H �V:E����k�Mm�F��1\��h/PA���{UwP�� ��1���o�Z�L[��]�i(S���K(6E�g�$���z���,
����h�,�sږ"�8ɧ�K�	���&�#~�ʦ?��0MAT�a�g��c8U�pA����:��Mk�	X����-����9�Y��Kr���Z9Ȭ|Y���!e�sB�=�l������1��=�qA���-�bj}�,�C|�;��H9
��%r=�|~�Wr����׸�bo�ZИ-��O:����T`�7$'T�D|��O=m{',#�x`�P���B�oݞ	UK�K>�Nk��M�p�qf�iY���faqvd�6K��#�eg�`���aV�b%�`3�<�����}P�����x�%�P�;�\�	8�v�0��p<�,��{�R{8o�>���'ܥGPȄ�:jIޤk{�]e�͐I��L@ CF(���p���A�1;��e緮�P�����!s���ic׌?�[�?
�Z(��0<�m �)��c��s�7���.�{��`]K�(��A�2��h�@��Թ�=�NMu���T-~���D̗��a�:B��V(�
15V�Ͽ�r`t�n+˝��4zrP^Aэ��đ�N1c���ӻ�6!�#�>o�BT:'(W_�(1JA�7�V��o5�'d�~tfz�3�~I�XaG�'�}\sZ)tz�"2�(���ޡN��9n��i1t [ޗ�كd��q�1�DQ۠�8�nK�p)8���
���X�5�GC0��i��bpN�m�dN�����y�%�9U&�A�w��a��u#�@[E����k^�~�u�m����J�l�*�e/N\���Z��7�M��j�A�z,���%%NBj�YĶ��n�&Yw\��KE'�L��OT
C�(2e[�I�?P��S�1s�>X��b@�Aǭƒ�Z��(�θ��X�Uv4�^��o�e�T׶�W	HlX��~�)�4�Z������NX�Ƀ�&�5�a3�ή�}g���@�$�Z5ٕ�8]5t�*И:�Ϭ���W�)�6��u�	�ex�� �`HO�T+��}�D/ӯ�\����BX��?�K�X-?�Y�m�C��|Z�/O���8��,>�d�%�}!>c^�Pk$����β51<*�4��%�Nf���q��ZL�+ư3R}C:jG��kPj��6�dM��̢��kw��da�lk�4<�w����CT�T�%'�׃�F=F�#�����vs5mo����R15�@���۞�I�?u�X^ �I�Pi�����ȸ��{���zZ�B�qM`lf������Z%���]>�`�ٟ��2��f���z��~��z�F���hR6o[������*A�-�Ywۨ��Q�qJ�H7)`܃�D��c�I���� �{Э˜h���Q��8\xB)2	u	�k�fU.0gl#���C:�˾:Dˮ/ц��+���7����	�@vc�3�P*JZ$0x[�6�9b��'�^���wG���lvp��t�|��`\��oi��4+�V0%J� �]�F����N�#�¬-�oW�G�J)���U2v�1��c��>#i�����V��1`?�iǞ���Wz���Op���	=5�
8��]ɊWo0��e�>�ͦVoc�P���C�t��z�S�j��S��^F�.��q�	�C��@�Ϸ{���c$9,ao�YiDڄٗ"*��C�*L�u��ㅍ�8�F ���l���1���O�'�I���u�u�e���N��2A�a �FJ�=�~������@=A�R���`�!�W���E�*�b�`���p��$��>w`ܰ*������x��1<�2|�'�<!ٝ��B՝rR�R^�cG|��#�!�!u|ѠDX����H�f�x�Q#ɠ��c��551`b����͚H�BC^w�'fĵI?Wm�"�'%�	��E(�ގ	����<�7�$���z���F)��Ma�?	�=�F�2��0&
a���9H�r�rS����}��Ič q�B(/��i�~~�جת4>����;�~�wT�u���|T�U��U>�����.���G%Y�����T���4&Q��!�%/�o�ѭ;.lޗ�k��8�q�$�	��z��Β0"!B�߇��x�>!&��v��X<W�;%��N�-CKs#&S��	���3ۑ&?4�sv�SGq�a�6ԋ���U+z_ A�m�����8ݶd��K�
��i�^X�D |S�)$��aJMx����88��Ս� n"ҡ�Qۍ�i���lFp!�K��v�ܓ��˖�kxX}tQ{�`Lݗ�y����6�`���U9�a��Vq��P���s�q
{� 5Qx�7P���Ӂ�Z���S6%S��%/i/�_���h�f8}Ji
�Q��ORfT,ja�_&wT!���p��}	���z�ո��to����XKƏ;j,k�����n��K�{�5	������6=��VFGơ�B�c��ڋͯ���&�b.D��h*���q���3xp��8�L�"߷0�WJbўi
V��̜:t��{�v��bQ�cJ�%�zSt9���K�,b�a�Tn��O�'��+�;�~���3�09�"�h��y��2�y���CK�o�p׶�$/	�Qa�I(?�������0kk��*���A���ř��l�T���3����_<�jODܱ�ٞ�*�;}d��B.�l��z����t�O pz�&f���`���-�߮�md�j"g6߾n�0�7� b�<��<'�}W���Uh�� �r=eV6����f�nڤ�3���)¯"�e�8H^��(��Ĺ�V5z:�f�%�S�g���3�Z�\����������[%n)s!���+�[=:Uxb����Y��N�|�ʇ�x�Quta~���}z�l��IQO,��+6�Ig�SƗ�a�[s���`Ớ���<��2�Mn`AS�Eě#hE�ƻ����JcL��~�����!��we��b"M������>(��ו,^+��+_-/g<�\��fs
��|id��C��_����n0�"^Ejʵ
�V�l`�Mr1t�!S�unmν��t:��7}""u�_�ܓ�6�.����hd4�b+�ݝ��"��x��]x�ҮѢ-�����ݯݫk _�$&���N��"՚����b�]�^r�n4�՜+!{Yܾ̾r�ƻ��Z�	�eKg���F�B_w�bvi�� ����fn.L��Nb���H(�ޢiWYs�I۫��N�4����H'�T��8T�����p�k,�����7���������/���9r�B����r5? U�2?L�=�Z���PicH�x�������2�=P�s7<ƴ�Ѝ���@���{v��=s�f	�@8<�=�M8߿{�V�8��gy�ɬg��g���wg�#�Ɉ�~�ȳp�{��v�^t��7/Ex����R\�~W�M���k#c�m���=ٹ�mbtK�J#4{LP��K�z����g�g��wقh�Mf}n�Ɔ�P[��Hب��]Yb�: ����:T�$��D+�L)�;�6����P��v��V�E�-~���)��z���k��k��`-��S���=�� ���/%���F��20�$j�|ǵJ��u�\�Q\���1�j��mZ�4�aGU����\0�<�+��Z�E#\��RCr���K+�Sⓛ��n�����{��3�ld������b;���P!f��F�,8��ܸV2�#������IV�i	�G�wcD���^����C�C�:-���o�ٿ�@|ğmݺ��֦S`����d��A�l
�(���A��s��� ;�X��|Aٔ ��c�Q
���}84}�W>Oi>3f{C3��1�\��.�6煻f\�Zg�8�u{*�	�`��$���v6��Є��\�r/\�jņ�qz�FD�H,��S_}Ƒ��4��m�K6EF��CW�y�P_V4��[g�\�R(��B��/!:�3�k���<�E�]�&UF,�t��8o��}ǵ���s��
����T�-'M L!�޾4w�d[��3�^���P��m��K��Ǿ�6�]��[9�P����%u<����oL��<~Ձ1`�m�1�0�����baq����<�t��~�c��Q�`�dˉ�h9o�pP	E�V�4,��W�K�}-�*�q}�����I�dFQ������:���W�&�c)z��G�@�W[��?<��0�`�~$0��(�#]C�@S3A�(6� e�u�ւ���d?(��P����Z��Y.8��J�P�'7���r�+ҌJdtk�[�>��`��3��^R�'�ODt���?l�QҕaH��xN�y/�W������?��0|3�p��4h�>�F��f�Q��/A�4�T�+9��C�n��ȃ�A�腃��(�\�XG��1�Un{�_l��F�9k焌��yq��tJ�HP����C⫧�����.�*�H�H8*�9�V�K,�%7&902.j��+?�/�S�"×,
T�-���t^F2�j����2<��ȓ�y���1�뛨�y.tT����a��!W�)�$x��\5��{1j�0Ȧ�(�#����\;��XF�1��l���*�ikԛҜm)[-zL�0��o��'U2[����\.0"(����0ZZ6*T��~q	-�@��R�� �e������G��"14E>P���" CLzI�o��4���1��x�T�1�:�n=�ח�Avi{�h�gΟ[�;~C73X�̦�ȩM|1���]���~TE�bbH|��T�)�p5~4�}n�'Lञ��E�M['Kĭ��E�Ҵ�S�Wq[�g��)�7ыs��������-lVY�e�_gFd&	�3��]u��g��$`dx� ǛD��ݏ,:�����v-��˷4�|=��ۓ}\��he�D�7�Гm�:��c?Ø�^�;X�^"j��?7��$S����w�oc7��
��o�Z~��%�	{L����[���#))_7Vz](ϛ\�0�W� J"ƚ{�#e���}��S���g^n*͟K�^�"`LΤ��P��P.g��ɠ�<\���B�n}�� 0%P�hԷ�!mj�
ͨ��ހsA��%��J���6_��X����t��ZW��,F�;�I9;>	+�}=T6�� ���^�.�v�Z$�b�@5�ji�fP�}��h�����bnofd�k����:p���g�1(��T�tm��(UO�b�H�{:�I�#K���	����;�K][�PН�9t����0`�,)\��@�ș�xJL��=�[.vY�p�6#CR���_�<	�4\�d��Q����W4Ez�a��>Z�E�.�=�$Q.Jx'���Z�74(���.?�ͩ;y����_�!���HŞ����K�Y�C<�I��,q=��u��t3�f� I}���`�~`Gb��j.��"(���I�����<������НYc`.����jS�Dz)�*��!s#��ۣ�:��+����n��,�޷K��eH�	��f��2ط���S�6�q���9��$ӛ�?���&X��n�����i�>�U؜mޘ<<�9Jl_�Q�.P;�w� �h�g�Jq��}����۷J��d�����/A�������6*:�N`�XIMXk',�%�I��f�������X6�چ�u(��V�ß��V��{��H~�c�������X�G40��J J�}��
)(��/)	��������9}������Xg��D`N�˖V1ApDWan?Jr�P��}𰑡�8Σ����ݏ��[ve���>[LFhJ�牒���1K��Ƽ?��Nw	��3��e��0��ulo5�#�o')��5/���VQ`�<����1.ʢ�#_�����<��ص���G��5qK�13`��rH���t���$8�y�#���Н<�B:�oS��+x�/�òGq�����&L��|��Vq{6�t��l��� t%��T�u�T�ʙ��#�O"7��\� i���L!��J9�|mb�0�|N�nT���{�{Os��w8Pt�j���`B`$�E���;����� �N�t���h�ew����5���T�L��6� �g�؀�\�m��[�c��F���c���!m�,��e����a�.]�js��<R�� �'8/*G��L1HR�I�l 㺛�2�`�_a�F�Mhr|��hW�g�8�e�������<yM@���-~��RE�����o&�x���'3I�6��PB�V���D��*3���Y��{qtln���Ī"�9'P�y��IV�X���B8$����|�����C��K��w�4��Ѓ�nv��j���x�,S�F�k��M�(Ѷ�$����,�+�S��Ǣ��U��!;�ncXT�hߐ/q�L.t���gAͲH�o+�;�E� �%�Y]H\?����g��J�jX:�HlI#rv)�@�S���O�(�#)1�p���s��/���,˦XMC�T+�e'�����K�_�=�uM7�&c��k-��td���o�{��@a����{2�N�߀�����'�d+��O4�2�<�Q�_i��~��7/��Rs� �_E�	��s��)Uu(�W_0ЧR�f��}N	�)6���N�M�Iw�2�N�j�Ϯ�Eq��is��0T�݁�Q׵O��V`��f���(����;hH�L�ڈ�]@�0!���k���]ݷϯe�6Q(�� ��d^O&͐����5�1�	;Y�2u���\%�AB��^��P�~͠��Zڎ��}���yO�'��7TKH�
*��`'����z��(��ղP ��R��\Z�J:/z����Y���:���C9H�jh���A0����z�����gx6�ӆ]��PRR_�e�I���1��Iى��jփ5�{�R��`-���d�5fv�챫(�"R��!��
�[�����0&'�0,`D֠����EZғ%S�T�����L�V+c�1��j��[��t}�T6mj�Ȉ�A^ܧ 0��xo�/٨��Fvk@+-9���V�j���N�%ƤM�ع�/�IΤ�Q�d5`�*Hϰ�ԟ�lJ��IZ��M)��#+��x�a5�'��y:�A��e�N,*ϗ���ƞ�x"ח�� 9�v�n*�bw��x8��"�] ���G{2�h1tm�R�7�z��P�[Qݸ\17�_��xmr��AvGTZGp���� ���7_��G���V����@�>�?�nO�4?	�ٗ�;��w9i��>5���5��w��e�	�y.	q��{�q���m��!|���E�n3�L��I-��t�їi��ą��<L�}��� ȨZsbHΏ L��
`��X��3��㒇K�]M�\ӗ�ݒZ�V���<U��<MdIl�=O��H��Qx�|�V>n�U�d߅�p��w�4ש�h��=�qm׷���
?�{*�6;��9}X�
���.�%Gۜml�����I\��C�����Ú.?�΀G�1t,�Ϡzt�u�.*b�� )v��"���^��:-u��n�9��G��� ��j6�^�zŝE:����pMȧ��e��[C�>�9�1����*�w�li)�O�E�G]��R��.w��#K�)�0a�/�8�$&��[\l�;6j���a�o7� ����<��!�᥮������em�N�ǦXD��Qa�eT�߸�pߴ@'�����؎��r�'�f�'��56�\#����m�KC��7�GO��57^����(k�4�}Q`%%��I��D��5f��>bm�	v���!��GASh�>�i���pc�{L]+�w��qszʖ��C��V��Y`_Y=&��J"*����ɭd�"&���r����j;����7�9���ߕ�>�D��nLJ�Rv�a���HE2,��u���|��p�E��h3�nM�Yu
�r���U��ZD����U]�i�~Hז(�d�)���'�3�;���z�kg��#l�mI%����R�/�(@P���Η�Sp��MsC%7S`�T�y��~:� �I��>[��2Հ���?�Ct�x��4�������Tr����g�S:���>�*���qm�[g�,=4�S��R���[���?�&���%
}��M��굘^(���A�oM��t��HY�2�0����^�%ҚA���q�C/�;�g��A>F���R�AG>�m���n�i�a�Y��똊�|)��my+�;���,+{/5��wp��I`e4��w)�%�Dn7��8�x�V��!��y��a�!F?k���]e��wfkm���#��T����=N�'����!�ʯ�� /8m[��oh��-s2��b�'�"������d r�"��Sc�U�'��(����Z|T@���O�
����i���m'�^�1�g&Np2�����(颱L��e��9���I`����c�� R>��H����A����d�f������W��u�D䶛�'3[5���v^����X�^�k(m�ZQ�!��p-��iƌ||�b��Z�̗�|�2��I��Z�cN�h��ح~���@�%a(09 f7%�9���Q:���K���A-����l�侩��>?��S�w��	��X��r�|?\	ܛ#ZU(��~��oca�};:���m�&�5�bC�,
D%��\E����C﮻Q��wb����|:��G�J�&xB7�iA����4a��Cpڌ`c#��߮4ʚ.��9^8$\�ō�+�#��@7^���P~䀭�ŭR2�P��ϒE(�fb0��V������� .���@���ϛ��>��r<cQ	�-B��_��E3L��7�=����	���5�3������{Ej�oR����������AP�����5�\�1|��\wZ�s�
ˣ(sf9,��"
u�Tk������K_u� q��q���u6�q�ƅp���RL<���4-�1��9*��T�C<j h_����#Xؠ[D���,�����%�ǚ.a�����_���s�9�8:5Q�1�-AemLQ��"p�v��B����j������,È!{�RY+Z �$��⚶��o�I�(S0�DW��E��8�(�%���C��M	�e���*��e��J�66yj.�Ĥ�J�II���������-��ƛ_x*nݸ*/�V ���`-W�+.��I���an:��L<�e�;���>���$߮�"*�#�?�g��/͟��g�t�@.P�Дy�Z٬������B��j�$/�X8��t�ƤQ�h�cl�s�Ʃ}��W+K��=�	9��[�W^D+��J�+ѵx��U�w��ARu�1�`�9淧��L���Ѡ��Em�N�3�����8{��w���w*cl<�(�X�ii�}O� `U���+����L�rT1GI�����[qa��i֛+݅=��
W��K�����
���:�����
�ٛNC�\��Fg*g���?D]W���H�t����S��ͨ´R��Ә��m�Y��-ף�� ���~|�K��չ����w�����q���U�ӄ�'}��*��Rp�:�
�1�:�6���ōоXI���Tk����*�r  $�y���)dR_t��l|�7M�0R-�[����XFF-������+��ov�����1o-�+s�C{$vu���O/��mJ\b��P�¤@��p�qx��T���}��;�o�B�\��*"�9Q�8�K��%Tr�Zɉً���[�#1�.n��1���@�6���K��X��{DL]] ;���uZ�Z-�t١vO����&�p-	V1��^$��>5G/tҼ"`L�C/2�<-��/�_�1���7q����;�avO �Z�>ꌎ�F9h���<D�:�Ǧ+��襆�4h����:�*0�Y��+;�u$q�C]M�����&Z�O@�O�8�ྰ���z�*o���L��5pޏ�tcڕ�8eT�� ����@;sz�e��fW��9�SM�u���:�F��'���e��b���jh�Fd K5gcI��2��8���I��_����3t�h�pV�֛B<�+U�K'����ٚ�k9Fl�bH�n��t�b�I�!�Y��Q:J�2O`Fv�#.���SѨ^6z��ȾPp��VM�8lG���'��t��Y�~��s�T~�1�=}��գ,3!��h��]���ᑙ4�������8xJ\��y������|�y�z=���p0�)�%4��ƙ���`�;�L��.���ܨ:K�߶�֛Y�cG�����SGwk呐u�)���ۖ�.ƆVYC\����y�J�Ø�4VH�̢b,����sa�oT)sk��V��G0SO���C-[�q29�Y�Qr�\b	� {��v�����r�(�Cq����,쉇�n�>f��O�O6>(�dHh-�Eήʣc�V��`/!�r[��0�[z��:�����% '<%�A	B��@�����}�gD�P_���?�����RHWo��	��2�M�X1Zgv�]! k���5��wba���9�p� ��{��T]zذB��/�//�R�$-%�ț�f�K�~��'���y�K&���9���8������
 ��_Ă0In�6�����e0�+u���h�[5ԁ�� ��X,p<<�(�����r��d�ߨn���7��!5i�62�Su�)��	�3��3���%��Juϊ>�>��M���W�eP�ť2���:�������+��X����Z�/Mv����4U]Q�R=L�נ��f��&��V���&
������e�W�P"@!�acu+%/	�N:V\��S��D�c
��fV�s�i/��چ�� }5��ީ)T�f �L �}�����'��E�M�`��)��&�b=����O|�F(�~���b,5�@�r+�~A���Jσ�M�^Y,�"��)�i��lU?D(�a ؀�hd�M*�P��[1�F�>iY��sf�g&�7��=v�×J�*��s��Y&�&�����~_��Wې�np������[���f�ҡ��\P��2��2mg�9.�Ƭ_D
���>p�&f�������4��|�څ����Z�vv��f&Q1j4%69��M��3����C��@��c��� ��P"��J����~��8��<P���a�)�hF���h� �i#N�5D[�)�wI�쁅=o�t��(cv'Vm�����N�t�C�G���?'%�o�:h�l��� 2��IJ���r�jd4�4Iɻߩ�XfaB��?�����bl��<�$u��G�D�$w?��Lj�n�Ӟ�:��"˹�D�ޓLլ���E�4���ܠ�M�`}c?�>9��X=�ȁ��3����3���S�k��?��u�PQ�-����lT1lRږ�h��G9�����%�Q�k��&����Cset��,ǆ�\p�+pj���S^@=�jz�Q�(�|Hݜ�d�-�gYO���Aqe[
R�[۾P�(�,  ~~^�-S�<�5aQk��
$�gѨ���!�W=�31��&*�vz���b�ܮ~����}�����ʯR+H��h~S-@ $�f��{B0~���=J���	1��u��@)� �̝`8�Õ�i��^N��Mm3��Ĵ;�*�ds��^K)��;����`C3U^d`��i�Tx3���\=N��9?b���M��f�j�L}�>U'�hg���F;�Q�c�ZO���6֏�x>�jz�G{�D��A@�t�g�`�F~�Y�H`!�G�����Fɑ�F��l�莯���"�M����UG{��7�tz��N��ᱬ�����Q {�L"�ۚH���(�Q�e�޹�G�aqÿ�ov���+��g�1 ���T%�S��r�z�;����Z�g��4�v~r��U�y���'�zG�,#�D2�_5Qgѩ�����J=pB���^$������A���Ic�-7�˳����'�8����ts�X��a�}��a���I�'.[���c��%��؁��p6ây��/Q2h�]�|T��q]f�M�MCr���k��͝d�;D�������G�/�[`�����.zU���'���m:�j���$|,�iԤ��J��ě>@�����'��~��392�7v3S��|�9~;�.5��d�أ�MށAɊ.���B9�IIO�t��D!a��	0�r��=� ]�(D�5�����#}�	2���B.��4�o>`8>���� 8����q�Y��bzbg�	뜋��B
a��Z�����{�vX�J|t�:Jxxg�0-5��$�Ǌ�D�|��������Fl�.aڡY�	h�׫���u}b�ن+ͅ_'kͨCof'_�J�og��^\w�8���"�����W��t�,��ܗi�>�*&n#�H�ٸε"�_��U��kx5��������dGNn�	�����`Zg�Z�W��#s4U*�G�F����	�N�8ӵ9�I�2o��z�����!�g��G��dZ0��a��#�Y)�o�j_:O�.����H?v�ә�'F!�j���{}�R9����b���E'=�Ɨ�{N<�=��%��]����V�-�1CՖ� ���qfFo>X��x��!�5���:qFUD�!�� ��[�u�6����1t���o�I%Ь6�`���p&O�;	�ьϠ}Kn�wʵt����AI�~"aT%���0�w����1�R��'���gQ����maoYh�A�ʬ�����.��}���CKd�A�K��`vE���}�a�W�C�zn6-Y��itr���ɓ�͂y����7�N�~�D�)~����\��@�kz�P1���$Y����v�Ոy�yMa����w��^1��ȏ���I8+�7�@�'p@X�'�*b�7��z'b� �ﹳ^7#��SF��&u������Q�O]��	3���h�NN坯l��N!\�eq�WFR4�h����O�g�I�M�r3��������K���q�RI gٷJh;;��=�RF�N�S6
s��,\ؤ��vu��d��ƭ\�KpuG=�H�p��"�õ>$m�A����r=�UŻU/t^�_~|G�$ȥ����f&[ B�(5T١Z	���V�B7-�n%а'b��W�|Uz�@B#p��27�q��8֔-l����5�K�������S�"���Nh<"���n@N���.9�N��r��9�E� R,�`�6u#5u�vwLU��-�2b�ؖ�� �\��i�٩����JH���i<^��&�bM��TO��~D�,��Z&9I�n�s�3�I��&�z�	s���j �00K�-V��6��0x�މ�
� 7�J�Ɂ����#����ޘ-��}����}<q����S΅�A�a�j�0�S��h���%>?,ɓ("ڝ=�y�K�3#q��z0�xeUf2���?s�b6ʉ9��p#4�@G�Ji�^Ҵ텨=������Z�����rE���!���/#��ki��&�={�ObP��S�|E#alRv�@k�
�a�� S�<�(\ű�����"�&[0�"|	05��̫��A?�'q�)����`dn�V�U��U�����H�٨�UlKӱK�V<��g�f���N�2�W1h{��h|Y��k��YUA�[����M{���=^��9og�9G��v�8����ڂ���P���0��%'��ۍe7?i]��$�����]zw6�ì8�4hn543�Fw�����N�p���!�Ƌ��'�.Aq����B׈�Y�&�tu���X��=�;��w���h�Lc �ͷ�,~h3�ݝ���� `�)lw�F�-�u����-��@\~fE�_FU�{��g�{�l_�E����F��?�>O���9�ESrؙ'�؁� �x^>�y?oM���]��M�����{���$�f��/K�fi���*D�"�'��[r������"�����������q&i���s�B~H^�s	��ra�f��z��%�v�V��1L�i#�Q�~���Y��+K&�-0��Z�����ky4�Fp�h�	�
�.�[��
k���C�k�x�˱����ӹsu��ǐ��=*i�']C\�3Y�F�v������#�V�TX/�[^R>���~s|��{�ob6�1m&0��X�x�#�EJd\ ��FǄ�����[:e���������}�͵��ހϻZ�"p�����Q�廥WC�� �3k�6)u��T2��MO�[GGm"���0�Bx�~^񸅽�y;+z9ؑ$3/h���]�����h���a����5��/>�����oUf�q�)��B��E��v�m��u._�`�m��րuL2%8��aǸ|����+�[bŰ�翲�X��n5�<߰����Ԝ^��OKv�`R��Yї�|�:U�;�$�Oƾ�%�?��|" ��-Fp���<���d�Wr	�G��b}�a,����IX���6`T#�[{a�x���ڭx�<���,�h���%LK���2���f�V���	֜�"���&�?��/���'1���k�o 	
�y~��1)��Zs����J,y˸S�=�~�N= ��Oz�� D����_�������r�`%2 ��곘I�&���݅jNNډ������`�q����L-�?8����bZx�v����E��X��و&(�+���U��q����[U��$�B���x1^�,�	�X����?�>*��7b7QBvѷ�=�s-2؛�Ml�v�"b� ^��,��5�����Hži�.m�y�ZZ�fy�=[��ڹs�A�W��)3�<���Ź�^�X�����L?�א����Z��?��l��b/n�s=��mO�f���h`�C�}(}f��1���*֔Y+ʡ�ꄑ�)檎����T�|̎o&W�g{�6�8|)O�0��Ke�  ��024	k�d�	��%����a�tP�<�e$�E�,��AH�m�C�]��Ĩ�-�Ot$�	�����-!�v��x��r:ˎƃ\�Fn�ΈJ��܀R�Sx �6ҍ/:�q=S����.= ����\/�'�j`�2�]��olp��swi�<����"�)}.X����v��\����"T��-;u]�C�o��C��"DU&Ε����{��0���2T� �j��Q�q��~�g`A&��E������/�x�ܐ-�0�����)�� T �n/ͷ��pO�Í�m/��vz��l��"�ړ9|[|��t��r���5�B��<C^q<A�{[52X���`��R`i�n+��7Mķ���0�2-c�x�; �3\���Wz��W��n}��'�<Y�ݫ;�K��M2�o8�.L���l��R��\�"������t;j� %n4�!�OZ�&n�,m�[�;�x$�P��D{���m�&��p�b<�+�tփϧI/�vi�p�S^A6�V�Vß!�)�Ճ���C�x?����b�Q�E��-6�&w���_K.{�G:{S�z�{�0OQ'2���y��$^~j��&J�?Ӷ��L� S �B[�>�M�\���ǅ��5���-�x ��!��3�)F�^��qXV��
��dYѸo�08~�0k7/M�	�b��zu�!͂O��¨	���6���7
�D��		��d�ڄ�z��������;F��<��1����S��k�_Ƚrb��)�1U����GA[��������9�Y�V褖і��`/�]V=&��H�����g��Jf�[alݙ�=��s��HY��|6���ʭ��J"�;����I��YK��Ӄ#zڻoq8�	���;����!������h�����_=��A1Q��P������% �?<.U��f��"j��%`^�23�l�ȱ Ct���Q�N��{�L����m��|�NIy�)�ܽ ����2S���}��1���Sd��G�OE���i�j����2�2�m���uL(���P\>l4��Y��.Z�e�a��i矩g���Y8��Zv��^�|1�Ĕ�B��������d�Vl9(��w�JR�#�eJFz���Z�q�%� ���i�U�ۀ��[?C�JnH�M�e�7+`���i>�L���E��
���	�1�)�8}TX���\��Ѫ�r�5�fA��Oy,3�UPx����ة�|xA�B�c����qIo{�C�bQ��YX�5Z�yC��3sF�	NY�5Ҋ|�$����H_'�9���,%?�e�,d��]!���ٵ��e�#�� �r����żZ�2%���E�zA״������~Rg4�BXj��R�	5(���g������^��� �x��X2��}.���H���:e\��e�2�YR,0:����G8|,-��΋hi@_�������)^���(�+�ON���p�0�s5��^z	�щif�6�u/����Dho t�k}I���ݢ�N�%(P7Y����aҚ-�����0�=e7S�/��{3��������t�u�R_�, �&��/_���@�wt66<�w�]��t���S��{Ӽuc�5�p�MeK
1�W��\�(&5���S��P��6-nV~��S3���^E��߀�T�|E¶�|��4��U��} ��|K��a��a��:��7o�	ل�kf�����6���P����P�Yb�l�1�p�H�x���$�h���=&4xI)�X4�� ��j�G����I	7��{z�+�Y4�-f�ۻ-C�'���ǉC��R�
C	)/���%	U��తA�ɢ}WٚvԢ1ױ���hi���D��1�  ���f%�$P�0<��SEּQ�����W��a�wIiN�����L�VEe�����J&a�`���C�E�w��ʁW.���e�X�2rJz�$/��VF�����~@�poIK�S�7����ر?}V#�.+�a�4hY:�-`�C�u��m��p��;��3vޮ�|�zA3�ռm���%0X�bY�?�+aYJ8�" fF%��k���O��֜��-$�����';���V�P�/��罧��@�(����W�֮����p\a����l˷+М�&<��G��>�*��Fp������\�N%�5�6i�{F|D9�T�E�A3�:�Nk�L�CmKvK�j;���1�1�j�a�慏���I�a�y�.�������l�DF�ICq����G��H$����J� ��D�z6g��b�5g�#���]�ﮯ�[;��㜍�gz���C��<��5��ޖʥѲ��EV;��C��3>Y�Ctk����!M������Ws�B��5Q)�Ml��
l9@���U3�`����<yN?J������M�(�Lz�0+)�
[�+���VAJ�)����I�F�bPBb�t��\�#y�<�����QPA؟ޚ�V]�?����<�C���"A&�����`P�/���jt	�^HpE8t�K=��ַǶv%9�,�K+-���"��z�	�*$��+n�]pQ��8WhUy �;H?�
w�j����1W�EZ��|��O���^<O���|�P��c�$i=���H���Sy�!�S�C?Q�i��Xm'$�_ۢ�}�w������u�@�U�.�=`I$ �����D#ͭC����Ho!���2��@��Pj��u3����	�M�R����*vg��I���j��+|;4��7��ve	�ʄx�b����be����-��6���Zָ��"Ĳ�i\���H'd�n�h�e[g�?�Y��Ĥ�]9��_�]p�wc^�H_HiBbU�|X�b��.n�^98��_n���g��2?\g*��]o�|�ٸ�6G��|'p��0���i�ȭ��\�։GFϼ��p�BPv�T����*��;�L�@�*�>ƅ*��&�ծ�+_��\�ڗ៦�E;� �G����g*>�ݘ܏ZȒ���v���%K���A����@�L�w�%�;ܸ���T�6��VƸ�";��ߜ���V��o��w�ܹ�D� w,0	3��Z�跂R,9�X�Ǒ6Ꮸ�=����h81�J�L�f�'�J�6��Mo?��iC��ҙ=O�{�1U�	�[��y��I�0�^%�H���4����w6՛����X�l�
��]qF$:"h'��^��g�ض���E9�e�݄�>�B�Vh
<.�����q�X�ۍ��Ug+�	��6&@�XJ�'�x�Ӝ$v��\��o둗�9g�-����4K'�wO [@$론�\'�4�À��p1�}����f�S�XA��L�܁퓄r����BOr��7yɲH��$���?�T斉�5�6��f������&�,\�p�����'XK���a������:#Z�9���	k?*����l���c�Q"e��.�6=P?R[bl̩apm�E@hj|4d&C�F���g{�5�M1��U��֮_P�I�,��̑{΁�f�����5���	�3?~��ξ$�_�81���fg�]2��X�\_1��6�յW� xVF���ё�f[�����	�S��܋N۶�?dx��|�V��1*Prc_]ܻ�?��Gd"w��R�"觃�7K��m�K�?�#�.�������a#Czqn�|�ꂴp�e���lL�/�!�@4�C�2�b{�L��y��I�ȃZ`,L�!�}iz��7ݡ�J��HjS���c
��k�X@	PgZ�2�q�(��q�t�g�Y�q� m:xC[W�1ߪ�_:��^��/I�t��+iT�:�b�Y\�](ª���8篥�0*�k���Dc�!i�>z3�+�x'�yC{�.�����{�G�����)F*U�s��ˆR#=d�P�<=��Ӎ��qeO�b�]�@Xܵ���/��e��!��T��Ny�G�D)��NT��X��ڸ�������f>���YhR�����aJU���Ȃ��.=m4	U2��͂���h��R�Y�-�1� WuVga-U2t\�3����/g�������c�@׉���wO7�p��N��7ߑ°�U��n�Z���p���bMn�B���J��K�t.E��}�zϥS���f����7���T|��C��0V������խ��2Q���;�
�ۦ�Oq�YT[B�q��4H��^<`�
�?�+aںL�F���c|R�$g�T'��5� �b��U!��4ڗ�S�X[Kɾ�/Q����8g�f�T3���,��}-�3�@���~�P�;܆`o�
ž�Ϡ^!ԛ=>����	,p�T�vi\vt��B'�kW,� nO6a�]>$,��0�܇?؂��lc�"���y	&��dmi=0������J�SH�E�T?��/��X�6�Sy�R]秭���HJI:{]�w��w���� f�8��fnc�^��ر\�X�7zY?�6��)ݞ��SR}Hk'j������5Q�y�̅�	�
�:�/��b���	�����^7��R��pn�rx�Sq4q��n�Ԋt?��Zä>�PW�	�[�[	��Q�qKM�W � �P�:�[�B��"����/�
��4�������I�&�K���_i=�Z���SJ�V�wP1����ik$+>��wҼ[�94 Ҷ8h	�|�n��-��%lO��s���~��BF
gK<7��xO	5T�	U9�;�d����C��?;�oC����|�t�����-����qo<g<���LE=��������F�5
��N�Q�6��`F���d�RW��֋n;�9�7)\Nm�Y���R�z�^?^�p쬋ϴ� ��U�AO��&�9˫�S��:U`�(����olJG]U�r0����Y<<��yb�~�S�u
v���6�3`����F����B�du86�p��nݪPB��L�Qm�j����G�{�N`����"H�6k�IbE�"ڻՐ��-�|�0F����e���u�q#�αQ,�ؒHq(��c�!�n�8�����QF&�b����1Afd��S�����SF���)ݴ�Si[u�x�SE8(D�.%W��ǜ}�ܳ�D4�f,��?w��Y����YLP��fE�T���PV@�ø�t�:�Ssv_\q�dQ�foJ?p�FrB�8�a��:�u2���'�/W��o3K(�Ɋ�?����.63�mζ��|��ws�����lyD����.����D�H��˳L=㐋j��t?��U��tZ4�;56W@4X�]�7K��a���>?���s��2E�&�Z�T+�0N��66H��µ��u�&����;�;���n�[Q}���L. �t�e=����&�Qf����itF �Ḅ���J}��x���$��awb�~>��AuM9�Wp�,�P��irj&8W��I)����� g�m���]c;�~+C��N:���\(�fG�d����F�Bڟ�mt���<p��*6G��F��Y�I4��3��Yo�I�3F����A���v�ϫ���I�F�A3T����8��]z�:�ZwdY���Yd����-�Z���o˴�f���O�ǿU9�ٱ*/��0�l��Ȅ\O��#�
p�u�_ON�?�sF���������؜��i)��F��l�"�8B�I��g?�Ч���%������CPY��o=9�^�{
�C�8��e� 3�u��ipz��d`��Bvw�~trL��l���R9����;N�W��o򧩇|Da��Vٰ*0�w�	ڽI3S�ꩥ�%���׸fl��v�o���f�4#=�Ɖd�j0UF�̘P(��
�������Uͯ:���豠^�$��3�l��c���ӏ�Kxw�I��(�-n����+MC[���^��f��Y���xu\�2���OH&@+^O��w�ˑ�)C?hV�Ke���3�o� �������UA~4w�ge|��&{��P!0f��Q��;��B��~�8y��$� �X��fko�OrPP�U�x��V����V{4E��iu�֖_�����d $�3���9�W�HO��h`j��p�H-�ڀ=nw�΁Ԡ��FN�3w[V9�o�*�jt�)!�`QEt�q��u���`攔B;l���
Wm�B�5�MZ]��&/�[��1��q��J$eaDG)�P5�ę�2$P��nu>'Йa�vQ��6,����r�#N�Im�R_�����=:��R�.�*���zhl��)O��V��$;�����[U5�3,eW���9��Z�3�C R���$�݁�>�|����oN4��������	*�5�2�Y�c��?uװ\}�R�b�|	���S�v���� �:V�Q�*�<�Dm����#鿏 �l�[?��Hn��qR���/U�.�����~�!�Ƃ�E.�1>�v<.���[iV��DS�?�7���&�����_G��Ml�>h���ˊ��9�/n�t�r^(<m���9ۜCwa3�,�HbC��k��F��1���Ct@�R3�f�џ�Џ�_���:w؅_}\6����7љ������F�"$a�O$�|�Jm�Q��1TvN=�}�N�[�%��EV\ ��Om@]v�!~/b�����$�q����ݩ�TLl~H�[��K��H1��D^�3��M��g^� ����,i��^� .���f�ae_3۷��� :��u+jh�0���5L�������A0�,b�E�x�����u�+�m��En�s2so�)�$�A^'*�T1<p^P <4��7fs�k�4�d�����tK���̣�D8a)�D�:�i�%ym1 ����[��PEY�)}���.t�?]�8��Q�ͱ�����j�\�j�䀂�,�2�&�Ea8��A>w�`���o�����w3{AE}��7k��a��l�	�<����m�Z5	 ���t���	�ѭ������7wf��
P��9�|*�h��6��B?�)cx�w*���q*��T6|��-w�8�ODhg_��%[��P&��Afx>K+G��.@δ�)2���h�6�9�Ex
�t���ln�p���nYS4:a����΢�5+�C���@k�����ll��CW���'���=�o9�+��\��w�(����9���̴�\��l7�[J���̿�B�:C�/���7�U����w*F��s0��L(��oSόh7m�����s5����f�*l
Ԝ߈�2����#v���V�;����~�^B_W���-R7Ӻ�Z:_��,��,�Q�T�{��!=�.�x��
�;>��Ƕ$�} ����a2&�`��Y�[۱��!�4�3��ˆSY���,?K�#�x�����/(�ыj�ʟ��5��u����}P����/�p�����1�,���������$�+o�
��e��;����B�!1��Eޯb���y*��6���]�怈Q���0_}l�2D���p�zF�롰��L���#�P��-6�Rv2#9TṮ�l<��Z���&ɮ@���D*T�,�qW1�kd]�'3�~ޣ��ϰ�թc����-c���x��&4�@C�|�������l��8�1)�.���p۱�&��|Q�%����M��9����j7{�i3��$Α[�-1��������[�ܐ�u�q,������{c�ӧ�T�=���#V Ռ�T-G�<k�)�$o\���Q��ڄ�:]�v�ј�Őzi7�S6%:`C2��!�ޯD�~�ޗ�W��lOb�ǂeD�`Ev����(TP}�b�>Vo����E����0�l�}�nPdq�nD�ˈ�P@�G�Q)���	p�N��mC�%���ə��e@�-�U�U���f�Q)eO_��n�=I��1��5�c��h|�ȭ�n����-��W��T|Ĳ����:��ːh?�����>��O[���.B���q�/R����cE OR��]?�3�"j��i)��z~R$/���Q�W�(lŷN`k�����G��Y�T<-@�m��d�ʗ\�u���)�=�[�1v@�9�x�ggϥ��tp�`5�UR���LʊXL�p���rr\������8j3dm?��[���#��2������0��άh^7��k�2?/ًaB!y�?Z�S�LCv�%tyyi���X�Z�]�W垕e� �bt��V��|���}^�J�3�b��^���F�Q���y���Ce,q���a���(�yb��ST���ج�����_W�!9�Q�K�^pTN2x���sqVC](��ʙ�l�ڄ�����Nt�����g��-��N6������M��̪Uu������ܿP�Y/�	[0��g�v�ԩ8_�P��"�o�ª�u��c�����#,�9���}�;�I���34e|����&Y �[�ɕ�X����ǪL���Y�\�kW$yi��'!3! V�
!]�G
�~Z(�r4|K�ۈ��d
������jK�tkn�����~J�*-������)@���綼���a�o՟����z����������;pK5׺�r��YF�Dꢾ-1v�P��!��_~�:�d���G���Ba��M1� F �,�A���M��|�#�K�)�`<��ǅM)^�.��g��l/v*�E��)uzË04�mG�M����B�yn�6���Y��d���n��Ctzo����+B�X�:6X�L�\[�7�rx���(`�GP���G�4�Q�<������Û2��	#�˽��'��k���
+�T{$�B�G�Ճf<�o��|���p���˰y�8f(�c$y��\.�˔ĥ^gufTN�UyJ��z��X��ݛ�X�9�LK���/s�K:�b��1��M�u����3��Ӯ��כw��"����(a�M���|�N�����s!՛�$�2���˓�BH]�"|���ԮDUÐ��O\ ^jOt���)�X��G�sa�Ւ����O���Vy�/R�l�!�Rt5�b"���=V{]*�$��13���aH�=H��N�M����~��7�O�Rf�8s�4;�P���pr����?S������0�4�˳=�|�+io؏�F&p�^O	GlP������%�&w�ݔ����4Ƚ�nϪ|�-�h� �:O3_���h0_"�UgV�i���F�T���gyK��iu(DҙU���w�[����69�Z#�|lX�W	|�?r�m�~�t^�,"-�Z�G���i��(�*�ً�};����,����o����ĸܡ Bq���9u�!��&ldၩ��>��Z��q�x[�M�9+�ީ�g�B~!����9��	z��5��|��sO��;�䁞�S���:U/�s�Xk��?���&���`�v�r����϶U@��J"R��E�b{�8C{I�i���Z�<�`��a�G��b���A��1̩U�_
�`%�᧽՜a�o�"V���eM �ø:��'U��DV���3;E��G	��u*X��l1w�i���$o� 51+Ƹ��!'ȑ$n�O�)�C˵�����k�́y�����0�$a\?��#3�[���+��M��{��]~]׬|b�y��ٴb�l]�UP�eC9
/r2�z3\��cl��� S͟����w���+5Y��f���������7wbQ�
����D�(u��H�F6a�rZOp�[������+b�Y�k�_@Nr�C�|	�(M��*���u?D�o�s�8c�t�I6�?�u��K���r���w}{)z)P��E�}��͖A~����0�VHk��_&M�Gn]2�6�ݓ&�'g��)-L�T�F/��%�k��7!g���}|M���=L�`zȪ3�A2�,�������4)��``t |��bE,-�՚|%	ˇ�*ad�(˔��y*͡�A*]_���t���g���Q���ʘ�˲��V��%�+��
��S��vR��J1,��ry+��\f!�8!� [�::-|��F%�/�k�J�؂��o��l�x���%M������=Ǝ?#������V��\pD��� >�J�*vN%$�M��BA�$]q�T⪴P�����{��1��e�s��Ìfp�/�W�wSr;ƴ���Ђ��t3M;�L��ce$j
=*�Ҕ��f����w�$O�}8��:Ʀ�O�LY���UT������hCh9�w-\��*��!*�&�RCS�2o�^O��H�h��O����lC]��$ρd(�ˁ�Hb��E�K����RG8 ��%��*=��Rsn:j	���O�\C�o
�5���Ӛ�E�����~A6ݐ�%Z>JYZ���C�L�_|��R����(�A�Ed�$�c��sR�9� ����N��#�0k��ח�*Jt{�{�.�iOZ�D�L�S���[��\ś[
dB�(��V ��I�.f�Tg7^��]3;��G�����\�N��E��:	Y׺_ߴ9j���bO��O.���b��2;�>k� }�N��yæ�/+@�G������d� õz �����{�8����<^	m6P���3〮�f��E �6,6u�-q�������sE�T��0�WY�rk$+FWQŤ��s�5�8 ���3d W��oR|��{\-��>:�}��풢����'��dab��-jq@����7��|�a��N���yy�Nl���7�bWC��pN~��ܭ6��nh�B�.K��=�¨c��.��^��fp����Lw�:D ]([i-W���~�E���CO����Wg��y-���$�矮�8vT}1�1��0@��T1���i��cD08F"����k@��������- ���WFX�Ara�C�ݺ����� +������t�>�Lɸ7�m�G"��O7_�l���YY��D4̋(���2�E�9������smI��\+-O�dz���H��F6'�I�	�6�2E���	�������li!j�S���J �)�~פ��z"7�Ѷ�M`���ț`��j�X�?5�Le� oe���n!�j�e-Q[&���bܵ�[*�lQM�.����r��T���}�;��\�:�ͨ�%�<���n�k~�/��3DZY|��厥]���,/��5NC5���v5�~���*S��<���1P�CT�X�گ��G���^�l���垿��⽳U�dO���vҚ�L��g��рZf���ߠ�Ph�P�KJ�c��b�-FɁ�o*k��MEm+��Æq��{�Ɛ�p��`���`�]N�����ϔ��
I��g��#�xe8$���RY�*Z<�đ�4��G��	/Y��dy[��ܼwL�� �'�% 9�C���V���y�?�6�pl��w!��V�w�U��X��Jn�*��(xhClX������z&0��i��ҒfW4��ub �����=��n�6�pc�\�]I��\ao�Ek45Ua�^�|��Մ����E�_A.��������%?�Ɵ2/�?z?C��8�i��)Ό��yW�AjI|��d�<�?C͘j4ku%��#�l�0��u���4����Ŵ�|n�wE(X�@��o�L�YV�M�դj���ss�3��[Q�^ή���,K9Zwn�
|�?& ��H٬bm�,�5�GF�����\���)ֵ�2w��N�*���
�BLXW�_�ˬ�#�j)k��G½�R����J�=� 	�?�ţ�&���|F�nx)Ci�|o���n��M�$j��qU�ԩ�h���$!lQb��	ݣ��>
f�6Gzd��uJ��VB�wմ���v��2���<��f�nL��oh^#��@WkCꙣaYc�ϔ�KrR�r9!�������z�H�B��?þ����+)�˽X�>ݗ�H��vX�����K�1iLS�K[