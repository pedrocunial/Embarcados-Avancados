��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c��u�KԎ���u�Ȑ�epih�+6s��+��J飁+r����h
��y���h��ܚk�l��^�t��ą=�-��OL�30�e�Y��Hsx+/�,�]�iUj\��w��: o��M�A��2ؑЕ�>z>�8P~�"�ݷD#���f�F�j���j�P�b��)��	6�omDz�N�ig��(j���(1,��������8H�{[d}�e�AA�=#�x2�J�$1*DB�/I �	&6��S���.�)��J̖�#*�3���_p�01��co�ݐ�L0���n쯈1�x��rѱ�T.�A��A��U�c'X�\�^�[��qx�{[8�$#v:0CH�XL�jLv�u���鵲�X��R����*g &#����A��-�sN�&U�S�Dk��7�%�
�ߢTǱ[�#���Ξ�΂���׌��]�!nߎy�	*_�(��c�v�
��u�Y���M�:�@��]M��[�H}���/��H��>��Y�b1�w������>��h�QG���v�=s��˜��Q7.b�����]����|QEJ¶�B~9�y���X4I|:�x�ePJq��ϊ��㬶�.���ǦT���<e�}x�=SoW1��K�o)��Hx)"Ffɝ���|�Tx��ɑ���8l-��<�?��G�1g�1�p�<S2�M�������F$Ţ�N`��i��o�"���ؘs�?~�Uf��r4Jp]Rt&9:�f[�1���pQ�FdMٺ̹���	��Q�n��@�RuT����hQ���C�_W#��5�x��o3�r�s�C����7�Bh r��e ?� S(J1�6A }ɬ�s�v�ض�<�]s����],)�&!Q��K��%[ ̱��"vJN���"Fp�X��kU��PT" 1K�4�U�&�:���¸��"���W�����g0�^_���!���$		_���ec5�ʁ�d�
i~�L|���@��	�WF9q���a&��Y�_�C�Ǟ+qr��gm$��|��s����qQ��¬)��lK�g��d��C����x�aF��^u��щA�'$��/��F�6���|�j�����,����?�˪��z��.G��B�jR�<�<-�0��3Mp�E܁�B|�L��У�J赗=A�4����"�Y��6�z*^o��|�^�2/[�vd��i'-�n��:�k�Y�7�2�6jY������(����V���p��}VZ��H�*��Y\��[�m'��y�#:�˖oYEI����3hl���vf��������qW��v��F=�T�ۡ��趀��	�|�y���(	,K�es�Q�tOO�9�uCH��*c�y��OJcڲ��5o�t�_�ؖ~�L�<@�|R��$NKlS�y��B���ڇD��Jd0���pya�3��H���~W1 �N�l}Ĝ����i��ﾢ���([��z�C�ȥ��z�$��C.E��ߔ@}r}&r#c��"�|�@āͻ�� ���k3|1�P>^y���p�F�Lj c [s#r��/�S���42ؔ�|?��"�λ���q�R:	��B\yq�1�<��Oa�DCw�Yg����:��ݾ$PTؾ�HG���v�������R�j��+���z�1�F�0�~�s�f �%�ɶ���}f�U��]	�Co������Ag)Ng��+��(x�F�F��	���U��~|H����)���Y�SR��/
���$����[h/l5Azے]�����c$}S��N�]"�<�y'\�n�Qg�c@��b��ە���ym�B��C�
������h���Yx�TEǡ>x-�vX��$c���Q�'E�j/��'g��Ő��f�F�^p{�F�b۹`I�q����m��������_���.ϴ���h8SX5������^,�n�W�٢��"0uV����3#
4���`����`$���jA����b �F�(�=d#<�����h��IX�/����H��[��[Xd��T���M=&D�}53�A��I=H��<�8�Q��{���>���ů O�q>�G�[��'����o��_N�.s��~��B���h�й����1��.���CˍP����K�E�rR�S��u��-��x�K�*�%_�NSQ<�^�$%2�NvC��6}u��Ç��T� ��ϩ|.���5g��!�a@�=2����&I wL�6�/�����E��?q�ɼY��9�3���G.�v��]��Q�n��i ��qvP�hS�0��#߽�{�ne�%)���4H�ߑ���� 2��,�C��27���!�+l[�hey���$����0�{�����Э�sH���#)�x��O�����T8����O�1���G�
��VR}�Ҥ{���(��nz��F�JJ���	9<>��ss<H�G���۴����雚ˢ�� ��E&QR��K�������=��s����6�E�����Ǥ(�p�V7�'%p,�M�۷Ɠq���d��Ɋ��zD6C�^�����;*nס�A]���~*B{$��B��8x |#iihZ͸��w[�9*kFnMZTZ<�1�j�IDŴOY��� S�#����d�̃���꾷�[˂?0f��,	K3�p���B�z}<g2 ��w<ha��o�Z�+��qq��<�El�M�l2��W�7N�=Wb׼�Ӡ�J�@�4G&��ȓ`�e��;��\s���䰟nƼt�������i�-4T��pk�	��Wj!����^}�������(��y�( 0��'�x&n'����V��JK��<Kj�|�nHU�<���D!X�*���Q�4dHt5��vZ�9[pqh���H���h�J�m�]�n�����&#��r�r�Q=�b�ln��ç�Ħ��UR���h�;�j@E�BP����Wuz#f��Z+$l�%D���,6��X�|-`6NE�n��`}�@oF�zc�a�;ڼM�L�̕�wd���2A�����ۅi�id����c�V�S������g����j����!�h�?�T��������2O��_ҹ��$7W�{��+!"Ӽ�X?pPB����	��ڹk�e�~��2��.�@�z�j'~d��'�h�MK�9�x��־׽RB��� F����P!Γ��5!:��.��oc��K�����3����=�xwn�Q���΋kخyEl=0X�,�n���ڶ�eA��0=C�I��]�]������N�=��as�B�}�hG@VZ��S'��Z��w�w���q��A������nr�}Ƙn�$���O�m>A����.�(�{
œ�?e�%��N����%�w?&A
{T+3#�%�y)�3������wn�L�V$H��b[5ߌ��p{)b���uk>��<m����@m�
�ݣ�P�D�d.��9�ʇ�!��;7�2�Ys=/�I{[[�O;o��K^��v�Zw�u�8�9��L!�`����!�[}p�8�;Y������{H�+�=-?Ĵ�}��%����L����Oc&�[��qŹ�����L�I��i��|�U�*(�|��ҿi�kcX	фG`�0��ń?SMנ���=��u������s�
yr}����{"u����JHBd�S�:VY�?�U?䷍�T���~��eHZ�m��J�b����&���Q�N�r�T�XP����🉙!��B4�9�~�ٗ�/�Dzv�����B��:�j%\�i_�����kx:�1�<7�5�h���`X��Э-s� �Q��vv{Y����q7��ϟ���nb2��B�l���-(3�a/b�[񡟇vE��"��T�o	����ݙ<��_g/d{C��gE��i}�z���P^a?[,�V��]7�.y���;CM��~]��oh���b ��ӫ̥"4�b�ة����q�6F�b����#�S�I�����^���'M���PD`BB�Ĺ��S/O$�����%:Nڢ�}�����YxVW��<SӺ��4�L�97���#�t_թ��\[qؔ �E�DB+���J�1��m������#ck�!X�,�!�ަ?x�}�tZ�ٯ2���j�	&���c�Җ� �j���3��Ig���t��%5�;Z�q�C�:PdT��?�Q}�HO�	�Ot��	C�4'm����ga:kI�i5s�g�ͦN�љ�9���恡����`,�����)�����(��x�#t�7�^0���n�
q8c)"�X��K��='�����+��{��p cbc<�=#M͞���@��!^#N�ԅ�Pc�C������7������:i��M)U㝧��qIv�����:�����4���v�-$�>�-�Mٺ���F�j")��|l(�[;$o)�څ���,��#0��(;�vO�Q6���VdY��燡"T�����.9���+[�y��1Yu?�\����g�;���d9C%�"�\G�&! �r�-丝�u�a�a&��0�A��rQ�a�C�������; Wq5*9r�$q���5�_��2��b��cm��폠�)�q8L'�V�p�z�q2"���/0�wBz/[�L��+sNs��O�c:N?��J��oA<)>�b�̻U�����ɞ���v��ҿ\"'��)����O��`�|Z�wW��ش�AHV�ǌ��)MƮ�����w����йD�
ew��q;�}��n����E�"��������&$�6d�����-����Dt�-���cM(��먤߻��gm����Y;����sڑq`8]:>�;�d\,�CtU�h1K��K�(ͨf�p%��ߴ�8Ϸ�o��(e�[��k	�ָ�4�נHc)ᜋ�L��AN��~m-�V����9`��:w�s5DUf O��-�C���;�n�M4*��	�:�)���q(�~_�M�@jO�R��pnsE��W�LAG����b����������)�h�0{sp��:/nC���Up��#F�<�����;� *��b�cU��Yo��3�LP���Ҥ�	9��P�~K�tS�KL�D�V�M*�t�����Q�I	�ŠN�%Ξ��g��#F/6Ca�۰���CbQ��D
�����w~"Ό�'�)���f�x���)����}�W9�hl��S�a5����u����~�t՜J0����0���ٌ'�E2�V��ʖ̔�0��L�U͉w4���;�H�O�}�vd��������e����K,&t��Mw-��r�hhB�hJX�ʼ=R�N*��!����%ux����|V@
؞V�rs�#Dg���������`Ȇ�<
�D� �-^9u:v�)N�=���o�#�8[Q�۞i�|GR��-�8�aa���A�ݎ�>��DY�e�'n˃%��$�49��������*.��(��m!�E��:/�]��������#����7��?p����bU�s��4j�ML��#�F���7�X�?�MJR���tMqp�U�D��Vf��������������Yݡ�*.cq{��8F^>ST�@�����������k�˰�.�hV�ʊ��I��S�p�0?�y1�_n��f��B�������S.��^;��ǆL�3��:�E�*�z) [e��F(%(� E�{�3V`���o�_�]�ڱF1��+S�`���4c�S�7k[�|���p^�W��p wD��R>���|L����m���R:l��c(AB�͚d�@��),��(al�����4&�������8� �X۷�R�^��t ����^<L�y	!:��c�4 ��LZy�G���F�*~�x��KrOzj�ܖ�,��+�,t�b���s���tP�.+lݲ�p|o%@Au{X �'��Y�/?Y��8�Ѳ�� �� �[OJ����ONS��AX��D.s�Fyʜ�?��y��� P��l���[(�Moz#�`�>3���^×7���ޡ\2 v�sm�I�I�#��_��:���x.��B���U^��#0*>�^������I�]�Ό�u��g���l���F9�_U�4f���Dv���'�v����V�����������F�5��g�"y��K��h�����`�F��_��q>,���/��,G��٫=n���|�c��%ڂ���V�7�c�6�����j�2���x�d�=9!Wn��˖C�ґ��A1���!q��.Y���}'k$�b���J�{j�F�%Hߓ���4�$/�����P�D-u�����&�����-v��=J�Lk�.�
�Rq��#�������P��Q��ľdx�I��ù�g*�.�* �(�9�k���Y�`�/�U���y*����z���
~
�� ��]%pPpI�b ��+2�A5�tj㪦a/�G��u���uL�{��S�к��	�.t�m�G+�V�{=,[z�� 60W���}O�ߏx�ˊd�I)���U�+ ���.�۴��?��A(L�z����J��x�y�QgB�a�=��ld�n���1��u�/^2�M,[�h��:D;@@e�E�OH��N��mk��v��
N�!��-Kx����Zk*dP��k��"��U�E�o����
}�)]d�=��s�W��D�',kd6�سD���v'���p��vb��"�AW�X1��`ǵF!����S��>�Cz�D�i��,̃���M�W6�	����:;�'�}�%`��B-3<Y�[Ԡ���6����^�BKWp)Z�d��_k.b��*7�	�B�[:�r5�����$�)���[1N�����Ӝx9;% �Ӝ���-4��Jw܈eoC=����������N���R"5H��3�q/�
T�o���s.o;�4)&�T�>�̔�����[�5	�������<�=k�RM·B���N��J��@���(��z�um�� z��=E�x�]�/�xLJ�R�Ef��ES���:�%�oI�X�+S��e�)���# �-ػ��(sƤ��j"�J�U�ap
�9+J����m�'@�;ZW���yX�Y�X�� ?9,!�42�n�u.��aq|��`��$w�?�k���Jc�63���[n��T�c�5�60�bl�ަ;�#��̨Mb����Ꜩ׸��0��݈�E��\�q���������܏�H
%C�}0s%��V��W�\��D��S��'���O��\	�jd��A�*��q;��;J�8gM'ފ�����E�����f�S�4��)d@'�'.�������-Y����-��gO\=:�)9f�Z��^���ڷ�"ѕ�6h��ӂ϶)��a ��}e�V�8�o6�9F�����b�͐��7�p�7����M�����3%��Iq��pJ'Yk�In3�laQj΁�����Wmnl�����KN� ���EƝX_���iV����S���į�ے�Pf��>]k���H_Qh�9i��&��?$����By�:����,���YH��{�U�p
�⊕�K{E�v��v0N̩wQZ�w�<)V.�R��D���*`tC�Cl�ć��C�;�K�:ظ���{�b(�8;�^�d�v7S@�rv�4�ms�Eә���U�����9��x���6-TzŬv�Z�1�ZU&��繠ض(�B��ꆃz|2�g����t��>6FN�v/]e��Ч�5�㟄�Ń��6P=�g�/2L�A}�_�b�Jm�`���Y1�	�����p��s�Xic��IF��V\����Tx͔Y��?JP��IyD�;��������FXlE�%9����N7D�	���GH��ez)�'��5�JXՐ��^��k/�;��'�L�\J� 1F�^s=�?�K���w���Ş̸Zp�y�Tiì��#����������J��Yn���6}���K��{�p���׉�\)Ɗ&A�SFm9.8��s����jC]�˽�n�Gs�#��j�&uĭ	d����}~��,��������˕m�$?�UƷH_w��HF�E��L�=@-���L*��}].�P�]�
w�m;��Ow�a:9?\⠛nc$z%<�`�l��A�K���f(�(�1_�oN�t��d������r�SYb	�ܩ1S�E���TUB�ܯA�r��#f�A)ߝ�<ZQ��B���]Snl�1ܱw�]�gfV?����9,	Kv�c89��V7�'���J���_=��.�s����خ�U� A� ]#(���Xu����X>t��0B�wZ%�/�!ܰ�ǵV��;�Qn��8t��h1�$D޹�����!~��"���p����;��ﮇ�L���v��8�G��ry6���n��/��Q�?>�(}������t�æ�A}���Z�f^�:��&~l�<��R5͕�5;�� �u�&�����C��1�2Й�'v��U2�_4*�3P��8����62(Y�������)x�"��^� 7��JU��͡��պt�2���`*�:N_h�C���\��E��)ֵBZ$=�;�pg[*�8�3�I�KP����e�9�]^���	�(���0�S��v��O���ޗ����n��
ۻ{�e���g��}�HTH>�� eW�!(�34_�H.5I�����?�)�+Z�G��/f��-}��$�]�w���yr{���.���b]�a[]Q;��2��A�`˄�:=!���T�6p/q�7�_.�˰������g`�.ݑ�%w����޷R�I���K�_�!Jm���!�@T%����״�4��9D��Q�B#��q��Q�ﴬ�hkf372��~04��ۋ��ܫ�ne��D��H��뵜�V]�޹��o9�2���s6�������H�6&n��΃����A)�OP����Z� ���A.K�р��G�u�p��/����m����J��\�K].��=��#7|~�Ed�s���'�6J���������e.H��#��	/�9��ƣ#Z��ւ�$�{�t�"�Fd��h��-��X��xL�>�F��[mg�-����<�o�"/��雼Z�rPH�T� Zf��dM�r5�`�
!�3���1@��Y����q�&�n���:z<���|#�cP�`��e8ؖ|�U��ES���"�;�y�:��r�{��n�ҝ�Z�0NA�W��߯qL�V�6�"�[ꁡ�Jl�w�����T��PZG��e�Z�⛜N4�.��N�-V� �3t�ؽ�|�O�sl�榓�'䭯;�	>��H[��z�����m�
n׬���Tj��������ԨE�nS;=~z��,y��&̽햾銫���#���k6i�:��z�ſ���tT��jc��ڤ�S���i�y_]ĳ��� ��o�kv��꣫:�kD��ɞL�j�D���;T�^n���afçp�6��͛rnJWK�"t����52"~v�# �mP���,���T*��r.����y�H��T<�&N�b��֊Q�^r �R@J xs�i=rc� M]'�D�G����W��vڞ�.l�}�y#͕���h��	r{�?u���=�j��\-����!�q������Q��`a8	QC���䱶kh gW�O��R_JZ�╒*-�t籜;p%�@`��r�ȩ�I���G&�X��Z>'j���\AEM'�$H�<g���ON ���k�"���$�,���ǈ���z�b����VJ�������
��\�ȁ��!�	AXv��a�������r_ɉ�������ɉ<�X.��Wɖ���ٿ �*T�����mw<��Ae"���<�piܩ}ˀ��y:���U���f��!�+2��>#w��� ߘ*���
�y"p�W=��vd	�U	�;a�>�O��箊:��(B�lH4�z��/%̽X/&_Y؋Ћs%t�!`\N����]<�R{4��".�An^�<��o8-5�!�Vk�2v�DW+���v�L�ݝ&�tO�-�����JR�%F��ғ�H�Fh�^:�E�J��M��?���Wq���c �o�<���)�/�R��O��<Y�ц�Չ��(�c+s���z���	�����ڽ�n�>�vÌ��e�"e|��P©��D���)�,d	��	��1�D������ko��,/5av�+K�OvՒ�s��o:#�}�%I�%dg�]>�u�@����;F�^E�18���|���ɧ�_I����C=E�;���P(����>�Qh_;_����A�2����,B�D�-�[?���߽�N�� ��Y�i��)�m���0��?[�7�A��(DM�e��ms����T~af1�qOD��>
�v۪���Bj�t�}^��hX��#�4��ċ��w_d��a<�_Ŗ7R�k!�J��Ey�v�YSd��$N�aՐ���n,ܞ����YO�D�b�(�ߴ:Z�`Ǵ�zq��\΀sK$�r7ǝ�
��8AA
�p��$�A����4�-�Qfg�(���'���d��4���fy���Ӛ�AtZ|����v*��t��u�q�׋�vO]���.�=�ܪ�V�6�|H�L:�����	@����+*���m��hPJ��`�J����D
�{��K+?#ǎtTi�L�R��!M[�Wx!�+���k�JX������H��Ps9�w���2Y2��(ј!�Z�b���~��<��Bt4�<įݼl>���<Q@->5ѻZ�.�+���oW�)NS�3z3(��pG�����i0g|.���r�X?��o�^�};���Sk4��<r�:��<�q��U
�\�1LnM&�_��qZ�H�V������|ׯ��ט7[��(�.��Ă�Ǎ�C�ñ���G�k�Ӟ]�i���DɃV���xɵ���<h�A�K�[H�pE*��dM,-��3n��3G4�Q`�x��P<�K�B�qD����3[.� �܉h����J
��F�m ��0O����6l>x s�-��Kv��"I�s��g;�������� }�_)�X�ߨn긌�C�!夃�߶�&���Ґ��\6���*D�IZvy�c��k�Y@j�#��*��pЄ�λX�4����'	�	b3 V)��{(�a�7��&�:5=��ji��F���H�}&$5��̔�X�ҏ�O%��2_]$��O<nl���ۓ�oRN):�w��=�I5�w��+9[,�Rp6�#`���ב���n�=�hY�T������y<I���k�T�:[�����(JJ�;�iǢ|KZ�_��aߦ/wR�c��"OЬ�i�1|s@^��6Y.�if�o�6��䣱K��5R�Jlo(;��y9F��$/`�9M_{w)hO��Qݤ/���R�$������W?������G�.7��t�'�����91Ń��IG�|�J*����iМ�� 1��_Dht|�m��9c�N2ϰU�`i.Z� ��bK�Qк�&�xס+c�$�/1��� ���A���L��>�-���ڹ!βB��O��h��[(�	
�16��-!�Rnן� (�3<.7�|�	%�6�g�� Ώ0�����5GqX�x�T�Ѕ�jHd�9r"����_�u�p=��-XA7߱\o��Ge�v����f�	�lie`A𙊒Lc��)��K`}r����R���+,	�jdLY����),����IsG�������;~�s�S�O?d�z��Jy/!9��ѩ�g+ȁ����Т�i�j�X�|�RMR�t:lx/>�����ӲQ��jv�.�T����d�<V	G��U�����|:3y}�A8�����r��{0~�;?��r2�{�����ae�K�E��$ܶja��Zc��'v��2���eճ5�ڢ�lg�v��'��nٗ�E�w՝9��]�c�V��r[�#"��ٷ��f���F����ur<j0��l1�f�R��}L��e�i��**TK�
�`�f�M�E�=K�ɭ��LM�0*RX{���Ђ��1R������1� ��=�1���)�r�^Z����C3�?�4�M��ӥ���L��M8�fVU����}T{�BDE�BA������o����1e�*�6�ZW�w���"���q	F�;v^#b8��T��&��p7�X�X�$K"��_�am�2��s� I&��K�RF��*�H�B�-o�O�AB ����=S|e�U/U�:��>�r�9���^V:��<��M��@B#l�IX�J��u��L�2�Eǎ��AD��E��T�c���	�؋
�L���O!�@�rY��TÎl�|t��(�����M^5��
��IQ�8?R<`�g�<���	�d%��L��\�v�v�Y��W8������z57:F��%�;�)�2A���M��(+����G� ��U��L��UP�* Ř�ߓ�/ƝG\�Q5jц��7F���,�w���oGҙ+O�u����6m�����!�K��|�vϕ)CO��N��̪D~�6k��m8��>�%���.�5a�X�Ow�O�E	ń�8��Lv��/��֛��̚%��0�k^r��<�'2�=�Bx��K�-�N�$�7��oҬR�m�d��`[7J�5��&ٍ�N�zd��iҤ��/|-#���k�(�Ղb~~�D�ėb�
��C����c���6H^����1��^4d�e�~�q��x.���@%�R,���'[�΀�5�����T�TQߨ��X:��B�#���}���5D:e\9�*���/Q��r.x\�{�՜�>Y"��_F��KǶ���]��\���<��{+�,�F�Rs��e���K(�P
s"[T2��Vq�(�ɏ�f��]�OO�\�KW�Z��������7������t�.4��EϺ�a�U�e��D�cswۤ�e��Ю.SB�w2�m�lBM.:е�nt^j�<H��H��O:��"�V]ZS$��σ8�W]�;��Zт��Sk��cO�/M#�5%X>��5!��60b���ŗ�|K �k?̔ܵS��>;�@\�eFz�~�pmp8�Ę[����F���I��[��Ws�� G�3
�v�`�UèQ��/�|�4Cc�(�-�R?{"��>"���\���nW����8ə�ŏށ���}����ӽ�cCya�D�� ��lJ׾`AS�P`<��.P|\�՞� �q��~��P>�rᎹZ���KA��`�Xy�r�zb_�m)֤�����.�ҔR�����I�N�#�َ� (㖤�UXʻ�Ε�����d|�"I�a3)sߎ�)�d�ѳ=�O�[ᬙ�<޴���$D���R��z��K���-��S�����B6_4,��_O%��]�-h�x��	Y��Taz~�8Q\��bͻ�Y��h�R����0��u��M$�aC�]���hN��B�9�B�e��9���	�#�Z�d˲� Q�a��]Q庴��M�\��}���ag�	�6>���2�/5Nv�;�����~�З]����v ��@��'M �v��0a���r���-��}*�]�˶=��(+��v�1���ı]�9�[�&�b������%/��y�!H�}�<M,�X�M��0�B,HF-/�U�=x�%�3n���gb;�EoS��_f�M8��9g���+zےC�br�dV�	����X �\��^:�c��s0�$���UhJg�G��׷�gz��W�!�� �Ma-��/N����,J���,��rB<|x��Ti���d�9�of?�ݰ��C���ҧ��GLuFw%�8Z�4�	�%�$H|� 0�r4�t��ۂ�e!��i�͜�U����v��2���b�7��6+ώMɞk;�B�vw�0�3�[���T���r�]əds�]�NF�l'�<@����K��6���<D߾�����L x�,��H�V~d��ښ\��}�8��:5o5(���A�RD$鰡��]�_}r<گ�Ť�2����¬h��a�ʌ�3���Y?'Z����&:1M 3��-T�ɒ�������G3~�ț��*|�whn�����.QD�b�5�[�8mz �!I�=����D�#�V)���Z�t�	- �@4N3�;^DLg��jK\�V��d�f���Y������h��^"T�2�\�p��� �k&c�Qu$��(V�;������gk��T/�EZ�ɷ��Y�0*�z��R�L��&�J�n��|�h����j��4�P�'&���UƘ-����X�a��-4�R h���箘�3܂��¼�X�P9�Zf�UC���?Rs ]��H��d��׬����;o	N�c酾�����Jzߵ����&D(���(sz��W��KH��$l�:�=g�	�˭i0F#Z�?�C��=t"a��(v�[�� ۥ�,�88��БV��t'/8�b�19m��j�f8��_���8Nt��9���I{���DJb�	L�I~l����_�פ��_�Z=T�����Yx!g��zh2�F^Q`��ڡ=�'IG,z!�C�:h�Ʌ�J}��m�������avm�Jx�a�)Лa��(��Ʃ�R�@�����?3��N꩑̕�,�DY�PnO1ٔD��,hH��3SR��l�Z�;�*ɔ�� � �m���pr��0�ӹE�# ?�MKZ�<��)vͤ�[�ۊ�~AK�젮�z[���֮!h�(,���mޒ�>�������ψ��M��z��f"h�KaM\`��ꡯߣ(��ë��+0sn����Z��[��U+:?�^�c��K�����(0�����Z��	�`P�F�8'��K��<��j$�Vdlf�IISř�6�.�S�ԡ�+�S��Ʌ�4�+��HZzՁ"x,�ϕ�[i�������<����f����������K,�[���KB�z;k��=w�.����D����2�@v�!&�u���EӰ��Tb ������Y�_�܌��펗6g�sC( �i�<D0�Qy���=�\�P
�B؆/a�t��?_��aUY�C��w�S�ln��l�e~�z?�1H�Ym:��&i4����ɭ�Ú��y��Cb��y��qtJ�ׄ�grFҾU��6�7ލ�)�W�ݢ�[�" �!��9~U��兄���t !�z��KQ8���_��7�
[�"�R~S��v���c*�8��o�Up@>�g:�%�`�Z�s�NW��+����(e�:oe����xQ"K�&�4��ŋE�#�aIE�oPdN������gd�S��}96?��+�M4�mZr\�)\�ey�o��̄�	A��З���öE� ԧ۠�O��S֔P�[��+}��%µv���*�(��J�[��j�2�nS��V5�?��E<��{��v��m�~7��%
���Ԕ�RtT��0q��aP?~�#.��j��r4�>��d��i0� ���9��u|�Ճ�S��,U�ئ@��ꪸN�_omk@@��G��@�Z"���� ~z�AҦ�`�ET����\Ml����(���g�̗��WY�컽(�d$m5(���Y~����˔c-~>�4�-�D� �wO�����$�1��s�9�>�ݧ��RJ�{E]�ʻ^��eQs{陋�'�֩�k�!���6�}�Β�H'l+��gٖy������5���yBǶ��9+��.������
�]4/��a������Z� �D啳���A��Z�) =\�vB��а����{�C�vk�մ=nwX�W� *�n�,��,��ঽ�U�B�n8M��f:7U��kD������3k�d��=�Vh'�-�خ�Y��嘼��ij�C������41$�����	�� W���G�rw��4�o_�_%����1L���C`^dO������㲺С�Tk;�H
�-��[9Ʒ(�U,��n�q�:ޥ��TzanuH���_O9�hq��R6؎yVt�	�I�7SvXV�X�f+t�Uj��Q'�?�H������_Ɯg�" ���nm!��W�uV��I�=[m-qU˲c�% �����irl�_u�{���nܽ���=�@��ux��|$��z�t��촲�f�ɞt�E�����Y+�`���Wy�ΰ3C+���+�L}L���1��?����E�v��{��QC6eM�Y�VH���d%U&��B�D���9 �lU�>l����y擅
-�=�O�WT����x|B�.ː�;e�M���b�^c��a����Y��g��o���5ٌ�η�~���fd���)����z�Ӹ.[b�Pg,0b��C�%�'��]���,>C~1Ɔ>�P�aI��y~q"�q�%Y�d���UΑџbQɏā��YRF����^}��|4�L�
��s��W a��*�
w�.(��8�����#�:���gD�}���!���gL:	�4�'S�7��'_^��A�n �1��,v7͊Nb��/�u���%PD��.�*q�aX\��z+L�!bđ*��A8�!�D�����& gC^���Ұ�dX��'��z܁�-I��+� ��)5�:;��+3�MW��I,�%w�%s�����6�s����T��s�ۤi�1�(�6W]�D3�s +?s��#�*�Nm`�dD)�ҙ39�M�?�RJQP����)P�'�Sل3F��;�4���c����.r=q*7�h"p�MzPZ{�d�ĳ��JC�md��V��]��m���7Q�Tm�h�����QM�ڃ�I��Q&	[I7d��*���C|�Θ��r�m���G%�N]uK�3Sh`������ö���ѓ\���T#�|���_����z��{U�����BoiH������ �����#"@$�/Zj�O>�Gw��)�[�"|�q�O��ݵ�	zAy��oj|�!�N��{�"�0�j�0AZfǛf\�Y$n��T'[G�5�_ ����p�3ހ���թ�'8�YHR���Jz(���^6����$���iu0�`�˵v���<���Z����*@����%v�a)�b��	(�Fs�޻gQ�R�6b��B��Z�p�O�&��3�,�`k�Jw��Ԅ��W�T�@�
;� e'��sj�����찿ڴpR׋�*��tk��y��J����5A��=޸(��MN@�Ryk�g�|�|Y!����2�����$~h	u�����t�,JeD�w�T��8�E�U���*�5	J�Ve�ä�4��+��߻��⢿�C�}3���@נ���K�/N{j�R{	i[�T��.��.�D8C6�'�����7��PJf�0	�NSZ�I���YaJ��zC��}�c�9G�$X�=%�ۤjچ�U/wg���qy E��	�S��'��ݸ�a����5 �C��e$�"�T��A���=A@�!�vvM��ɿe��l��ͩ��h0���b��y��-E[b�����k���Qa�1}V�U.�B>��Y��q<���MEzY<;��Mp5,�$No��{/��������k�j�fR�F�����.����,T�E�sD�^!���^���"��C�(��������,���Ҫ*��~ B6s1��8���SJH,�+`�o���h0Y�}p�~��E|j��W�w��InB��)��գX��-����[���]M�0%e���A}P�I+Ũ��|QF���~���r���SS��k��p6TT���U�'~9a0�9E'N�$O|N�d_a!ց�*i�h^�ia�cj>t�ykck��p��d����R��>�*�h���2#E�+�������;��M8�$M��.!�U+['�>��N�au��ʹPm'��lu����~Aá�䃛;���J��{���&�F��U����\ݡOu����c֛vn�x�X� ���F�ΐ�����K�;�N��.UAl}Y�x��B���̦d˷�,�4C�a����q���
����"ݚ>����!��_���q!&�(�u�)@f�-��~ա}����8`�rX��>Vf�:�X�y�
��XD2St���I>�9��%r�R��T�z �P>4�����)<��.��~RF��!^5���!���A�ӹǶZZɴ*,2�@�_H��L���<&Q@sQ�Z��zdf\532"��v&8��l�Y�9�M�1Fr{���4[�$f������Ƈ"�T.fjPay4�Y;�+�5ܭ��� �S��DE�ʖ�R�^L�Er)�~���VQI�k�d��r_�UN�Y9G�K�;6�8�`8�S�j����Af��8�3LhSZ�e|U�n���C%X�G�F������оirm��j��?fp"ӛ���c�䕔d���eT��G����uBu
t��p�	)�b	���1g�$L4Q=���F]�����O�`|�߷�E}��i���L83�զZZj�CE:UW��=m�00g�4Q���IV�w�/�2�f���QM��Lj���Otd�����Ө V�L����q[�󠤼\dp�&s�!i�vP���ʝF+&����c=��rZ�?�c�;NH�TYz��w�MZ��E��S~��%c���8ne����y����&�<�u������EX�������(�"&9��ǦTR�3��|�����[Q��֡���}��+�y��Ca�Y�K��E?E����;���un���i���`�Y��	� ��
���Mz�8͆�m��
E�Ղ�6;䮏�p�5�圣�Η3Ҕ�&�q/��ן�]�P��{vN��l���#�jKw�5�RC9T[�O�������/�o�Gt�IM��C�b8YsO]KކH��x��.��� ��m����CI	6���<!@y��4�bn���_*aKۧ �W�BpiH�'|�?�8C���^�ﰂʳ�'���1���T������^�8[�R*i�o"�����* ���f���c��.����D{�^"��! W�ѯ�E���9jIB})��^����P5X
Mpm5���etA0������QYu6�ƈ���r�f��#.�vT|2��C͊[a}���tT���3���E�n�S#���qj��7��VK��b�hԳ���Q�06 (����Ţ�Wy������i�Ը�JЄ�C�Xzg�!i��Z�@�R�1�Kg�9�S3�ĖO<�giKh�8cES�&3��0��_��kg<�A^���ᮻ�m�����t��i��f���!�Z�E�M��R!�2��d�5�+/�-ruӾ`3�K;���#&���$W��[Xorу��>�'%�A����]�	G��sW�G2�?A�����t�~S���6���$�L��3iu��2�v�Ʀ�<��������]j�E6r�B���\.���<��y����\F����ݮ�j�C9&���BC��b�� 4�s�:��C[��[]*nJ�k���i�|MI��9�$��?����8<�DE���ׅ1�!M��`��G�
����C�.Q��^�r8�d�2O��e�蒣E#��B���wdM6��N���!�Z�{˗q���\E�Q)���<��6�`Y�Q3,I��+��+��|vZ�uT�(���H�)r5�y��$&���8y�i��#e�dP�/�S��a��_��0_�
J!�#�xC�`��ᶚ�Y��j'Eh7Avc�Z�/v��>�߲�ōݾ��D���|��O�A�w�����lb���,wB�w��<.�09k��x�ς8���$v�dF>%6�f�Ig�z��
w��?� ��W!Oܙ�;H0�5yWc���`�(#Kvf��ʄ����5ꎺ�8!1�Q����.)���W� Aː��,��߫��@̎�PLl�K�6ֺ��в
��ۑ��3"'Q�7�`f[�א��DWd���J�[�Aj�̇3����D��)a�
�e��u�n ���C�3�A~��[��Xl���E�����hq���q��O�@�&!�<���^$zy�.���@5�=!{[3����l`ث��i��z��)r%8��#��/\=k_�j\�d{53�����%�z�lo0;)�&X$��U9{����)Y��ul(|�fsL�B�ZW��E��һ�������u5q|�ȫ"�X�tM߂����&?%��v���%d��r�*��H�+KI�w��-I+'�'�=9��z���@O�|=)�qf�O��+,?Hj�}��!t�����gK�/�ؓ$��/x��%��x<�\�E�y����lp�H�8�k0���@}������5�uo/�mvm6,8�A����~SH����ԁ���'�+r�S��y��b˝n���.i�[��ܜg�E��s��#��r�β�(DE䈌�~����'���p�*��r�n�Dk�H�]�<�b��Id@ܦ�n�K�y[mhi�[3��n���gk}�&�Q_���1}�K��QG���,���,-�vS[d�!+;�`�� ��Ez�m>[^Zo��i�� {#N��$<x�4��v9���d�J�Ϝ���%"�����;{��(]�����I�<\�A���M���b�q�c���]�a�nHw4Q@�����m1�2����_�����s+�-���"@�o��s��ɧ��'.Mh}NE�+�I�)���K����+C���
Z���6·�V&�����Pu����c��\�3�	\x���@��[��P�ct�����xoԏYx�I ��d@��S�]�����N�\�S��VT\C�D���	�Ωh)"�7E��ZN���_Y\_>1��&v"g���Z`��
xװ���6 ��6����ۗ��'/��
�3L�9���,��%RW�Qx����}�ky��|g�j
�ۺ����܎����������6�^- 4�F+���9ͳg�ek#ff�4�^�	�^�Zመ����/�V[#{6�⎀#�1�o�@�dݤ��(��9� 1��e��_*>S�@�Gʠ�����ԉ?��k&���}�zb�p�>��) a
�]u	�o����T����5��9��d1e���g���f���*H���]T-�M?.����"!'⽙���>'�.����y��3�f��}7��I���<$�B�t�Ac"4�љC��T��X���L��0s�r�A���<���)��7�?�UA���ڨ��5yf��̩>�HwA����넗��j+J���H�6�,�bK��#�B���pB��'}��VH_�U2���~��r�0u��TF�p�\�U�g&�������edz�>�h���SD��	h�n���_��D����A .w���`�.���uwl2a^=�x	i�8B����&�O5��W��Th����;