��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[����������=�U���*!�;b���$��s�>ր�<B��щ�QЈ�8��7;s�gNE�lU$9��S�ڇ�F�K�ۦP:ym&e7����nt�$3^+�g /Lx�E�\'�l�ZmH��g��D����I)C�� a6��w�n�^!Z���,E�7ȧ���Q�;����4��&�CΗL5��M�?�V�qwi�zF+�qC�5?�vn��`'���otW��������ubg��D���KO��D*����z�z���tj��80v�bݲ��5CQŭ"���\�C�������(a��I������ѕ�V���/3g�+�Ҟ�����P<=h��٭i��9�J�/צ�c��v\{ck��Lc0s]Nl��]��\��x����Z��X����,psD����ς�Bc�E ,8p98����/~�~�"X'�n��sc\��3휲V�u,ؤC�C)� [���X�9lɾ���ҡ��{�ˣ�m�j%v-&$�(RVB.I��x\۪q�6����DvN�9��
��f��\�/�]��u����"}�f��"m��\S���k�����$b�!:T�lf73$h3�H�4eRk.ɂ�\B9�����5IQ6v�{ۑ_h��V�\MksOš�\|��S�[;��Գ�$΀y<ob]���Ry10[@�j)������Q��R�#��z���4����S�~2�j�ϵ0��%E`��S�`��A��>Yl-��׼-�6��@��쀿�'�8���(����-/��@j�p-�v�M4-#Td<���3��\y&P����k)�#�9i����#�c�W=c��Vp�#���@;A��	�k��o�m\]�����x�2ݕ��X;���q2��8H���#��FH}�r~�W��zK��ws�VXՆ�z�V���\�6�N��'��j����b*�H,�s��%06�繴�̆���@��;eo��M0���CX���^O�3��I7��O:H����!�m�O�r�j�x1�-�i�Fk�"���12i$?���.j_jTml:�/�`�4�>i<ꦭA\���rgZC�B���&�R�]���-�3&��MQd�ꂵQ+������j����5�fjӪ*ʓ��pu9�=��T��y�<Ͷ��Jz���߬�4x��� e8�]�B�	�8�?W!��U��ꗒq�>����c4 ��@^���F�r�È�sE/M%�k`���}��$i�5ue3�+�w9)�y�÷��q��դV�q�ςGBQ��ֶ���*���6�}�/@kS����j|��l�)��Ԁ��؞���+c�4qmR��8-\n1s ����QƖ,$�:/"cU�	�*1��
���l��HS��AJ�);��3�Q�Q,q�:����ٓw��A�h1�,3��:���|$��>��mT���nw���>���:��?�at�Q�#a�7=2:V����k@�$H������@E��2:����8x^�A��^��(*�W�7;y������d
�R��$���U=��R;�=�Z�&��(ӭT& j.M�����]�g)�,��?��Z�t��˸�f���	�AJ�N-7oL}�`a�*��#��ȏ!��禣�oy�ꑊ�4Z���-q�8H�����(�ׅ�,�(C��0�r��B���_���"|^��Iu�;���
ȵg����ލ�0x�' ���o\�v�HR����oI{?&��Ο�h�/��zP3GƨۿE'���=���?ß/���+x���'1�O9��غm�ki5ÿ̶�;�r�t&��-��FMK�/T��h(��(],ϱ��>�~p�<��NpL��(U#�s��eJ
e����ˬ�ggG�;�UA�qe�2�~4�L�$��]e'���.k���;<��D���7�f�(��Ao����	S0�2����i�X�稆��yU΍wU��`�ƨ���y��(�h�.eȦ�3-�����QvT"lϙ��UU,�1�Є3Dʁ���I.Cᆺ�)�+,�|�w����#��z޷�,���ݷƯ�D� #�,.���"b�f�ގ vt���:o6d}��ԉ��/.ݳ#�*"���`����m�Y@���!��1�G]m��5��:��|� ����`���X,u����e�t����ċ�b�8J�1��P�0@A�_����/���,������k])����q��^P��W�x��JqΎi�Af���w`]�0�uȅGW�8�>�c�� en��ڜ�.��:�c�pyO2b��* [i=�E���`�8?��ő +�R�4����<���Z���ܸ	=���}�ǽQ&�o�l�ߘ#,*��X1B+�cv])�A����*��4q]-X������$�r���)Yg�<�N�I�����~"����b���Dg�V��H�����{u��ib���֘M���, �/�0��D�2�],HŸmqy�(F[��:ަ�tű���Ɋ�N��Y+5����ak�� ��X|d2���e���|�no�VU��!��x��U\�5F+(�:�R�DCz�|�GA;�ͼ�ϰ}'�Â$�F��k�'�|nvTtov��3ӑ3	X��j��n�dX���&ī�—P��3�Lb��.����5����Z|˚c�ߒ��Y%<<g7�vg��#A;� vn`z���$6"f����|tei��{���>[��dz��n:̸�����5$���5����&��>�A����t0f)@ڛ^��#ŧ0ʺ�Q�Vѭ�UI�V��eP��VRi�/Ӌ~���p�o�NS)�����(�v0W)����$ �Z��t��Y�ã&�w��j0�@�Npa6�@�QL���S�T��N�}
��������m�Q��bΘ �[夤�bB���u{
���m����$��X�t�1�l)�\Ę���N��д��)QZ٫�^�ޕ~�MuI���J���<�ӦK��N���e������(�)���$�P�I�#dh*�,�i��p2��昪T��IyR����C_���|3�?4`�����.W�y{�ɀY ��!��Ud���j�b1Yv�3C?z��dPA�sc_魿��t3��K��!�L�A����N9~������/��m7g���?����c��<����,�����RUx��)e:{�#�mH*�I�\�^QP�f!s�v���@��hC�԰��i��t�/��~�����=��K�bi�\��g���=ٔzt�bRE�*�"ʧ�l��T��,�*#��Y�~��oZ�YAJ�ޟJ�rX�`*����	S�~U�>�jo��Ax*��E��m!����!�Y��Em���&B*5@�uQ���*�Q�_�Q � -��fY;�{5n�}�12S
gL;��L��xZ]γ9�k�`}5��`rx2��|�*)4���+a=3`������zít`3$�{�l(���.�9~"�+ ܷ�BJbu@�)�{�(�}�B��
	��\M���B����e�M�s�U�|(�"�(xG�ip6L��B\�ʄ����랟�֌�� �ef��zE���a�*
��fJ�2��L��x��>u���Trss'���?�BN���CV��݂=��K�S�S��p
�KS�����2��A��_;�kMR��C���~�/K�HV:�:�����QPpM��чL�9�F*�����n�s��!V�Ì�^.d�b�A.�	]��h����i����O/;ҍ�i���*��?�g��p`�0U�_aaD���`C)��W�# �џsv��W[�~ۅ�yJ��PU}��u������88lҙ���љ�2�;�GI�&���#:F���H�݀':+:�z��$Gp����J��{i�U1�UP��g�V��$H~�ѿ<;`�2s�J8?@g/Y#	P1�V�@W��e�	���,��b��&��,���4!58a�%�3P3���؄仔s'��A)=�,�F� ��Xe�bY��+��m��{�:�,%��M:�<���7k};�*`Ԑ�x�$�۞��/��~�u�D��ao�+4�B̆����]�r�PUB�;�#�8N����0��������z��ɸ�c�s3�G�iE5ϳ��֤� F�矺m��u���Сa���
��-oU���i1+Pgc
���9�5�a�"݀����W��V��7��iꂸ,>S��YtV0�ʒyG����W��lq�Q�j�i%�զ�����\}��;��̄�T�7τ]�aW���#�jI��[P��I�
�(���pq�k�K~~=z&D��(�"-�X>k�jU��G��g�	��_m��c��}T^�v�Ǥ�N15�饍���jf�Cp-I�
�������.sw�5S�g��7�_��(��7GR�O�I��Ӻ���3��j]ca����=GH�é�> �!9tzro�/��"��C�?,�㙉;Ni�H����d������r̵�}F�u�f��س[�}۝knx��=�s���й2���z$N2�Iq�~8ݥ�`��7����S\A~��ɶ��1Q�&B>����z��E2i�+V|-�N�+x�mP�M_��J�`$��k�X��M~�����δ�ᓃ��(�)M���7TN1+�+
�M���3�7�΅��(M(�Q�u��~��"ҞD_&���j�w}�ߋyj�C�1��HP28�s#��&���������n��#E1�qo��<��?���_ڌ�~�,�t{�Y���@��rEhvg�6����Z����_Z��p�co�mYTav�����^/f]�� �Y?��^\��+;9o�v��/C�X%1};}?a矬v��h�?����h���/S�z?{�}>�*��SE5�s�!Ds��D����Y��US�=�b>m[BF:�v:�䵏l"2���W��ū@ĺ�0��h�S��a&��7@	w#mM��Ҟ�mRtNm��Vz��P[ILޟPwd.7��D;{U�4�up��c$&U���������5�b<"�q��t#��-�8i�UbOl%,����Kic�C���=w�6%3O��x%⮃��~/O�H��HWG�C=���vd�v�b�4tJs������+&�$�ق��'����~�.��Ny�v8�UX�LQ������B��3,���%D����y�f7ҿ)��߬�M�D��"��~n=-�V#o"�Gt�q�vӠ4|Ү¾��_�J�߭ �t_�=?;[[��5�A��V�c��yER
H��\>�e;W�l:u\A�'R'�#��8.̅F�S�f���%�nPG	�D~Խ��O�S�il�f�|D.�����#eU���8��sn�G��%g��HFo8�>T��y{�K3�t��3>�|�ۏڭ�R���^���Wd�ZL7WWʗ-	����*��Ze9�:�¹-2
���C"EF��+ړ�	�k[t}����\���6P�ސ�{�5�hb�3�������<�K�����#��9.P#Z��R��*z�:�{���d�7�n�)&9�y,���F�=G�v�B�P�F���1#.^�+���]���]a"���$`�����n.8q���Y=ɸS��Ћ�&��f.�?ٚ��Xe�{��?�!�v
A>�k�RB}{��M���Yմ�d��������,�0�Td��z����� Yr�yj���������	����<:�?
��b���^�?P�a��F���Sf�*[[$��BΖ�]<��W�Z&��\�X*^D�F)`n�;0BZ����W�r�_j_C�J?�wd�ݯ�0��,�Ð�>c����]B��o�x+���Mm�FZ|	@?�r�ڗ���L�]�	�NՓt�(������7#�[�Z4�NX}`����X�=Cr�G6v�
�zI�A@�r�E�O%55���FlP&�����%F-r������c�D��hwËU0V!����y��C�Z(B�3>�LS2V�`u��Z(��0<�~-[��ɄN4<�����N�k��	��vAB}�hfi	�S�vb��ED&`{���ݜ-�
Fr�ˌ��� ��$F�la�g:9��xeW�)	��9�rY�P���x��u�{��Y��z��ݝ7[	˜+w���%R$�����a�Y��n���;j���ef:��A�x�b����~:���~S�ј>@^^�C�{��:!���ngp���MfOZ��ؒ���2���]1�dNj;�]~^b�ً�>�&�(��F��z�`v\�TMj0$ݵ�����}=��b�ķ��Z��gs"��N��Z^�DN�SMY�˫A�EW	�$��x�����YR&�y^d�9��I.	5�AҌ.��W:�њ��9��:,�}>�v�W��i�ۈ��7�*=i������(a�0��s�b�H�dơ��^�D���s��Ҩ�/q��V�Y�����wbmcb��|I��K�C7���G
(�pv�:1�X�n�Y:Fx�V7���H��G%aA��Cϕ����p�,��A�A�}*�u�k'�`B�2���X[@�	8��B��-2upҔ���*���4� `�_�T෻�&p�x`0� *�Y<�~��ua,�ՎW�8ɛ�2B�6�C�o�\`��}0s���e�o��9���G��>���8n�ugB�K�|Y�L�S} ��v�d ��['����

��k�Oq9�
�Xy��%������[rb��������9��O3��%����uM���B?_�?J�CKhJ����B(���E#�|��,Է�1�	�9���m`���fJB����v��:��W��!��9B�[����>8`ssy%���(��q=8�9�]��;89��?��t��O�e:|����)�V����%����y�eX��E�V�,�s��׮:D���p�	��Fa$���&��w��I��0�b���J�^���G3
�s�Ҷ	ɾP��
rMЦ�ʫ�Yw�4<c4�*� ���g�/v�?
o���?���K@�p��Lt[_�*Z_|1tY��t;��cH�on�{�e���'��Q/<��KR��l�S���rn������;��|r�[��-,k��ɣ1O
�e��)�@�뤚w_�"c�<�L(�@v��'�w_P��M(�ښd�K	�r��|�����j�Ƨ�8���������C��'y��,���!�K�;�̌S�Ů�B�)���.'�J��Q����k�6,i�ҙ�dZ+���k3%������F�բkG lH��}ɕЂefcl�@����;��� b��	����G�o�dߍ���PJN�y��7a�=Ǜ�	�A�;��˻�es��<��[�HN�8*Cu\���[���o�|lΤ�(��c�D`�K�k;P3���ʔ����@�jV��k��mp��R�H0J�P [��JM��f�{�����3 9�n��Es0d���v��.��f���*�$6��2���ņ���؂��	�y�wv�2�a�H�ާ3-��8�	�l�I'�4���o�}�r����	��W��Y�[HH��n`aU�7!5�1�y��Ț���
�aSţ�&$L,O�7D^t�V�=��4e$�ݠ{N��4V���7��~şz0��c~�K��3��z^YR]U�,�C����ͥGڇc�����e�bp���I�Ϻj�gub�`E),�^�Q<8��r�=��qJ�!:�h�+rg	S��1X8�LQ��nJ�Q�ZaU�0��6��ni��n�6�F?��D��KO�{�W=�]���ΫT��9�9I�!L�+\�oVJ"�ec��n��UW�u�Aꕚ�.X=���ed����-���6�1ap�q<����oN�Gz��|�L�eS�S��f`~��%r�N'L��i8ǯ��2���� ���>'��W፳�D�9��J��eTYëɺ����	r���)Z�@@>k�'
L�٪����R:���ܹ����ubiO�UԾTp�L. ���`Z�s����tN�U�P���6�<������dT����a-n���_%Y>�� 1ҷW��ٜ{�ҝIW�(�A��f��;6���%��n�U�C2���m�T�~n�`��W"A�v�I�0� �C�qTy�Fح�>̷�6Ӧg��ڌ��F$�
`�Up��gB�r�$���r���MG��2��ynU��݃���۷R���`�ˌ� ���1C<�q�t4��T�Y��`�����7�i�f��e@->Ɵ�����/T_�[��ܑ��
Yʐ��t�4���+�F���i�����%�h �y��d`t*���#��?!Pũ�B�]b��W��k�O�ѩ�y�S���p���(qQC0m�rcO����I;��U�����ڭH�F�ޭ���'����i�"y��,^$�^�;�P���YH3��PhT@g��D4�7h%�I9~#���ls�k�Ί�Z�����s���͸��A��V�� +,a�?�
=x�����z�v{O��=��1�ұ@F�WV���*�A����4�4�AHzq�ml�軰�sx�-2>�/�w'L���'k���3�`y�Sz��7�8`7Z��o߃}�ڣ�4%��I�黭�h����ދf��$m�uFqʇW��.�@�V�#T��kK���/q�����X�6{#$��]��.��oRmt>K�X���JMF �s\�B/?T���;�k�J��N�a�q*S���_���:ҷZ~��"�o�`	�KWkMU�7!�S�^���+�H�� x���m�]i�6�x�\P,Y����v2�z��a�%�"${F-��B��9�&*@�3�Q��3��0�D��h��/�`9�+lB�hX����m�r'G�tT�kd�9�*P(ę>����%.x�[�*�-�6 ]A��!��wp�����d�uv9��i
9�Zg�ޗb�L��+��դ��J����:�E��{��2��g]��
�����j]���{��S+�T匱٣�_�	����Y8Mt%=��0���\���Z�0������݃2�xY���?
Wn8c#��!�<(�5=� ����鍕���M��lp4�u�t�@�C^=܉���]J��G#�Nl|�r_���C���,�� �MS٢ڶ7�_��a&҈���=�N��:�k0"~\���D,	s�/�X��)�h퀚���`�E~Ts��3��3�C�J�����8kd�&���q�
0]Wu�s`�k҅��^m����>ƿ��S|����V��'G1b��ONV��]9N�HTi�`#'A|o���>.��P�wu�	���h���;���\�fN�n�q���~.�ĭ�ӝwU�p��E%T\ *�P���C}[�9�q C�O������Ф��]�;�N�t��)�)�&�h��?ݮ�L�B�۔.0�dn�^E>tB�E l�O�$�`+&'��D��%Y���\�NJH,#����)���c���}$z�v��?��עm�~*�KҜ��O姅랆�;�9�9���nP��K ���]GdhE ���Vh]��Ӏ~?��n�5��&���g��!r2��O�7_����g��~Q�/�J��@�Y�̸&�M4�e�o �r"�(/u0�g�r�KxQ�E-H�"ak�U{3���fВ�<\����^��ιu�,���I�n�}Z
�i�~�����I�p���O����и�g�����gF�c�Ԡ���w�P�{��Ɖ�������VhW����|�]=o%�^۾63�SYD$7}V�(�Tg�tB�6خ!R�P-uKa�f�B�{NcZ?>����wϗ��!����H̨�=3��~����K<���F��P���V�;�Y�g?1uM�c\"�@�!K��i$4�0y�����pc���6�翽nno���(��,����^��;�?{(�����'햊+B�~��i<՛ԧ(��`c�����~G>}�$'uF±�R/DG�~x>	6I�7��o�g����m<��q���%c�Q�R5���D���,�o��ǡ��>.(�1	!>����A�8؜�����_< 4�ӛ������S�!(ᝅ�IpШ�m���_
���Pcj�m7�-����G��"�M�?���2z���Ml��},dOP64�ĩS�3@��/�;�/<��xt���uUٹ��%����� 
is��j,�S���
�^�J��Rs�~%��#����5Q��7�e�HC���/�#̸����2��L:�dӱ�������������L3���c�ݻ׻�\�KGт��D���U8�;�<���M��*J��wO�Q�����O����SvW̍4���������k|qw���8�E4���>$vn�h��wS墽�����l��I�4й��蓇��Ti��o��`_j�44P�P��c$�Y^�@gW�>� ���(g�l.l�m�8�X�b�E=��WC��	-�[\��|�:�n� �'�Q��(YԠۛJ��@,�lgh�`$]�7U��o�Ċ���$�+�1rn�r����wm��,�$�
�����(K��hz��_��FK2i��i�O����֜&�?�� *��S]v�PB�7�R���ɚ��i8���C�4S���lEC�p˝&E���&k�=���s��	�v� p�.�8�b��w��ҕi7ئn�l��KB��.�����x�|\@(lI�4���٥�~,;�=<��n�M���(�k0ex�i�n�w�7 ��51d_�\ڡ��HS�	���aa)� eM�4��Y���DQ93a�� �Vh����g��f^��H9�9��y��=�o,	8w����#ջK*\>o*�Й����Jg���"p�;N��؛�gB�<U�w/V�[�;M�l�����A���+����M�]�I�a-�pf_[-J�ZtC�#_�'�	fk/�V�Y%�b�m���~W��"J�Ryg�s�l� ���4�h�13�C�G,�@`��ٗ���n�oM)� ���|� �ºHemXWE�>!x�caX_�ش�s�z��fX���k�o�K�9P[�T0�٣�y�#�3�FH!�D�#z9�u*��&���Hٯ��J�1\��v�.��4��{��l���c����WC�s�a%h�?�.q�gC$����8�B��X�5�����-\����N�._Э���ZS"k�h�6t�s�=?*-3�Qc|�o��~�F��ٱ&/�X�g1�)�1�M�ط`�v{GZc�˘��ư�_i����3�<~��9]�:qt�2��![�5��'/���O�̥�"���2Vq�a���f�m�z/���4���'����[�]N)� C&��LAW�F'�B:"O˞{�W�@�m /bN�v�_��3��X�k�a�L��>Pq���":�	\L?�� `g������)��v��f�?s�i>�_`T̻��(����%�=Y�ͫ���᝟�u��K�H�n"��O�o:`-����a��fU��f�,��w䘶8q����:������ם�ܝ�� �v,����ֳw�z�є��\P� �W���j�cx�S�mH~�j�u+���\D�Qop/����s�)��-B�����xU'M�D�9����ou0d��Q�P�sK4=�����)0e�+;5)z�/�S�F��`BA��F^�F����}Ƒ� a���M��sdrr#8���岢�m���^�d�ɍk�/�b�e3���kG&�Ŕ�._BX��+	3���Ԏ���߫�9�(g0�n}�	Z=P�.	�D���얍�͙�D*U�A!���ܮe�F��b�B�#�xOq�x9�x��M�f�SR��K��[f�q��
������[J���ERu�Y�4��)i�~1�"���쳽�e]�����KaB�|�ϙ�ǃ��W������{�Ұ\*��;�N��ϳ��H����b�&��c�$#��$���%�"��f_�,��ʓ�����p�U��e�|��+����)�q��<tV��8�mh�nR`D�d�:P�Nt�_F/_T��x
࿮��e�	���KH#���F6�Em+������o�GY���MkemY��Q��F��tAst]J���b�����>Ύl�`���l�bgF؜�HF��`ʄֲ]u}��Fc��Nա�����؝&�+Gu�t�W�`�H$����
J�t�C�`ݳ�8	�Í0��,#�E-ף�7���8�LG9�}�U�ΎVn��f��C�)s����R0�OT@oh������5�o�YH=Vs���\Шȁ���0��}�����ٲ��\e@��-GW�zk�q�B��MM�/+o�
��֌6��T��_2�e�q�D�m��~�_(��]3��ݺ���
�����3�����@�<Yf�~KO!�&��^�I����d<��`�G|>���%�Z۴�TY�;\5ڜ�����Eo�dn&�8�� ���y?gމ��u/�@�����$����f??Zg0&�a���M��N�s�&���G�Z�ƪ��l����ӹj-F�D�)Q6����B������I�pcC!=��<����a��ۧ�@:ŗ�Q\qГ?�F��4��L%x�XV��r ���Qz̼��P���3,����z�UB��ߟ�r�	�c��nG��8����Y���T�-ؙ�-��#�luQ��n�]�$Ȣu�	�r�%�6|��+��Ȅ�"F��a��M���z��/EǮA *��~��yR�I���#nt5�_�����I��ߧ�#�<b��P~j���j+�(!�iJ��N���w�s�e&Fp�CI,BCY<�!Z��������s!W�5]�\�e]���qO���I�Z�Z&��X���m���5
��C�;���S���H9,��7&FY�����)�YO�c��y;�����R�V_�}���rB�3\�6���1�吝����[�ઁc�U���L _ �H%�h�B�����6�7�[�S�����X<.�CB��n<���-RJ�;��"�o����a��~v(�K�����̧�o�
k=0X��mx�L�ҋ_�$R�f��r�yk�v~���j$ڦȕm�ޛ���5]M)ǜ?������t* pџ72���w�2�lȞ��h�:_��7��ڭ$Q�U��+�b��ES��"�C'Kb�8e0��ێ9�y-.�f�0��N���ȫΛ�1o5��guMr��
���H�Z��yZ�&�E��H�A���0��	�C�#�,d�/�9G!0Xz[KnUP�p�=�\c\V���:��Z��EJo���BM �<4����%�����4��,�H�Z�5J�DpWH��x!\�@0n_�H)m���<��k�|�te0�)��r�%Ʋ�':�sl�y)�tA���te]@�6}�'�?g�b����oH`���
���d6>����(��%7�Ch�O
����C5����8�Fˎ ��%tk.>��U�������:���-�m�úgbü�~��N�ids2T:;|�)L�Ha�m�,)4�dt�+"�o�7�2Xl���P������9���q��V���n��QvS�T���oOC��깮���,�~��@��i��>S���[��+�D/��S��KA�����${ab�\B�����D�edm�^��>
4��o �O�m�}�������1���3.N�/�m��O���Ԝ,�ə�w����]an�r�Sf�ȼ��i	f�/T�L_���5�Q���e�Qִ�˜�`�O^�p� GZ�|�z�lt�]��匿Y��/'���S�i����M^�5�������3yF��0�����
`�C�#*^�W�B�x͟�.�g�M�=��	�d"|�g��L,RZH�lomş�E�砾�<߄k�$=/�3�6M(���2��|����c�\:N��l1�'�Z�"�w���⩯� )��6��^ǔ�J��+? ��|T����"2��{�[��6n�e
:$l�rﴽ�xh�`"$&�v�42�b�c�;�D W0�h�豁�*�#]kH�i�O�2A�Qv{ǑЭ��@|4+��۾�����s��x�ݏln$&}�}q��k��*�ݽ	TG[�IU��ɰ]=����@���3N���i��]�Oڐ�ͷu��
Q95M\j�lS��UE-�`�,��I&z�h����^	N.�+hJ����^)�ܽ�+ޕT��z���Q�wK�0\���=����^�2���@�T��`DI�Q!t[�}�� �B�hlu�R�cӰ)����,����d��{hXlXA�\4������� �<�
x�`�'x���O05�*>|�V~�5EsP���ǳ��8�?=�Z�F����|?�ŋ���v:����	1P����x�s�������䶓']��&���^�"��g��6��WZ��
�<�m���ͤ�4Sa��z����=�E5�))qs���@����,2ù�f�?� �Qj)����S����4���:����%�i���لR<`5f����,��őL���z�;\cf��k�V�+Ũgx��� Q�oP1eP�+���il����#�-���o�_���6����:�-c��)��g���{sm�j5d��Q�y�Y>~wo�S�9�G���,�g��ơ���@��J���~
�R��Ȟ�Y�fb���-3����՚]���W��)��d�B���aM>�j�P�{��r�旕HE����V��1���
�oG|<I�9	+�\�����)Uw���r��dTL�7��,�Ln�� v6�a�����V+ �&xámC#����Iʊ;��x�?
*��c��	�ݛv0��@_N�~Sd���� *בs]5�s�+*	8�`qA�E�\��0F� ���?���%�~y����[���k�̡Z�C��@�A��F$�j����-W�κ�	J�~��>I�D�Q�D�O���6�(�d̤N��+3�df'�#t=���38̏��P�x��?���+[�����(4u*m� �ӿ��U�U\���99����ٖ�;�mߛ�x`��D��$ĬL��{�ԭ|��Tt�Wv���f�^�4Ӭ^�͝L���y$�Oo+�N{�ʙ��d�i�\|rE|3�V�'P��5�݋)�����S����5�$�{<�j�U>,+�U9�<�����S���L��9��j��f�ҟ�ؐx�W�)��à����/mĝH���{���hK����L�>}k��ب�3�ILdiLE�,��nC��r9���Dn߼�p	rي��.+�lJLf�y���c�QhP��s�������cꕪ񊋿����G�hcY�9�
�L���T�,ü8�`mY*_��<y�{-%V�#o]�T��CGQ���R�4�G��/��d������!ô J4��᭬	ջ��X[ؼ3?�5R�rY|��^{��4r�-�w!���#ַm;�3��=�<,�6Ϸ �`4� p_k2)Exjݒl0�?��&���L)��щ�Cb�D=n��V�I~
�~�]�0�.�sf��<�)����8 nY�h�����y[�E-�qW�R�a}�rW����q�|�]�������&I�ө[�ms=�rkݪ�T1;����&�� ݢ�ٲϬo�ǥ��X���A��o�}��|�g��t�������U�N�$��30\����p ���H�Wm�߷����07]g�x�P�k	�.�b8b gHW.M�F�V�Mi�?�5����ÍA��ç[���'��X`��rV�va��M?Nf�;ef�^��D
H$�M)�v�a�������
`�Pg�ތGT�nQV��;z��S�sW_p����`Dt���k0�!ғo�9(B�$��23�gP�o��������wb�"�_.���,�x��m�B�J@�$��������=��1W���EBܮH{�{=��f�Eь�	x1�m��;V���i/���"/��`�`��&d|����+�+3�3��9��_�`!�*��/p���s���ds��)^�s8c��CX���C��ϳ��vb�$IS���5�:*�=��3����ʒٮ�[�<����|LC���[���������:�QҶ��A3NA��IG��W|����e��N@�0	m�(�t쉞4kC)��LۗF���	޻�׬D���}o�	F�b�� ~�&��'�swMW\e����e�ƻ/��;�Fq��@j��yw7��#�+�dw6�̆{`����~zEڿ��Oa;4�h	�!����oeJ���N&�w�T��0"|��\q��������s�G��y��-UxS?0 y���|D%a�7
ͺMw��eIN_ܨ�SVW�b��*����-�E��.ŕ�l9Bi�pL�3D;��c��V:�A�ҸbN���h�u
"f�5)��\<�t�P���3b��\�MLɀ</)4!��!��ɼ�g��`HpǶ��ӹ,4�4��/v���=�9X8E�����&���������x��E�w�<�鶶-��
��Z;<��V��_�%  �BmAr�Q^�k���w68T��J�/^DB���Y��0� ��>�e��WLO�o��&�Ń;�,CFo���Cq�w�!��b�6j�Ә�k~)�m�Ӟ�Y8.���k��),C�.'�Xl��|��rlo�Ɔt���a�x��1��g�����(.f�t���oB�=��6���K)����;e������BH����("5�a������D��--���9%v��Zb�"H��M��։ ���i����h�Q���%m:cJI�A��0U�u�\�0qn8���2c�%P��eq�Fw��-���`��e/R8�h��υ��Y��"ث-TS^\�n>G��p`�JR�:N%u�<h_��ʊ��8���D0�XF>���p/�vt��ÏN"7b8����
��,Ir�{�('�	�C�3� ��u1}}�R��+h��D̷s(/�׌A*$&�Ռu��j�Ha�kXq�̺������u�N��y�]���K<��BBmZ��m�n�L73ѳ3�h(z08kp�&-�e6�����:o	�a_�'g7�m���J��iW�=��#mU���ǘ��u�6�;�0�1���Gc��X��pdX'4��ï�c��(�/���M�/�,�Ol4�i��Bt9�~l�V�w�m)d��gp�֝��||�wT���5�%^6�{�G��𮏴+�q���X��Jjy&U}�	��-�������@��ĕ(��J���m���@yf	2�̓B��:�\��gK\E~5;�����)1$yڝ�O���D��Xv��e����o]�1������#1�A�#�o\b�.�J#��-wW��r���������,�v3ہ��r0�Z�@�)���,�Ss�$��V����_��ez���g�^��9��k�L�"F��u���(��h��,J���A}�H3�������V뵽9*5jE�ZS�'&N�M��C�8n�?�mנ�������\��v����ݺ�L߾�h���m뿤~cD/�!�R�9���~��s+n��޳��
���0[g�Lߎ��/����	j���)��^ka��:n�5�+�#�҄�'�3�� J����EpPF�R<߇Q�TM���󯈀-�D�U��!�@�|�;�K��C�Q�Ծ�s�GaAKYhRS�٢�� �ɾ�ҙB���
y�g^^D����I����#=1�(�"�eu��t�B:��,Fin�9)d�����r7���>k�lP	��H/���S��i8�5����I�(/3��̻��)#6��w�.�ճ�K���'&G�).�?�Չ�Nӕ�b���h4A�(��1D�в�ch�p�|��M 	5��ؓ�㿥r���� ����K�c9w��$�i�a�IN�<�q\hXL����B�1\&4C������!D�6b '������27�P�^D`D�s�ps�ZG���*�Y��B�����"�m���K�=�Ou&�t0A��P����c+��㆟�2���B��>���&�uGi��M��X���߲qg]/r��7>Ddʉ��$��oO����\R���֝��ܞp,�6Gj0�NmM�'���8&�
'^�	�w���ξ�f�QA�`p��� ",@��c�5ʘ3�a��d�<xCk���O�{Eח&�e_�}(m;C�4�Å��[f�ۻo(�����`ɇ�^3N�+qEn��+�J��M���YW�5���-7����*U+��!�T���ˠ������#|�,	p�KR��>�3��H�S�&��|��F�d�el���q3H��Ca�}��o�E��m�,�0������1��m>h�Z��M�M�vH �V4	^�7a��1�N#�
�V�n�]vT�������=4?�M��<��<֒Qc>l����K��[L)L�Ul=� E�,���������/�ow�˲���tE{d�Z�Nln^
�	�x�[n61	�;���� Ҩ��w�B����#���2�����r�|~F��="�6����Sfd�ھ�����K��j�]̓�[!�J��x�p���f��&7x�līji��	�i�܌n���,4z�C?4�K.�B���OQ0B5i�͒FU���뺤�t	��K�hc���q�[����n�n�q���3Y�T��X �;pH`�N�k�PB�n5�5�sqqha�Lr{`�2��/�Z�9��+�Vi�5)h��?k�o3���0���Mi5)q�ɔT�L}���"��͗�Ib� �A�2��bo޹�ۥ�0�	��X�����Aw� ��U��z� X�3��V��i��0u�j~�T��>A�O�M�+"$�V��~�P�W���}����B?��ɾw�?0�ˈ��*�G^&�}`k���%?F.�h���r��$����v���]�4��v�;Q��W�!��$Wec�7� "���-yw'�+5���'P�e�9�D#��-W�8�m���������R��8�'��g�����ȟ��P�0k����$�)"��"�{�A8�r 8��)�)K��ұ!�]�e�~wc�����P����L�/�<�;����~�A���{�1P�x���X�8��{�t&-���1�w>�/���OUߔ���I�ј��ݤ���߇��*o�$����' 	�T����vbT砈p.Z\�Z�oY����\��Y��tt6HfZ�Ψ���گ&H�|.�	�����)c���*��:�A�{(^�%C�n�_��U����:�˵h����8:��j.X43I���n5�'�խ��1�d��)w��^�DHS�"�V`�?
��L�&�g)'ɴf�N�e���J�YB�V/�ٸm0�a�X����޹b7v4���<����@�r���Ou<j~pS�3�?ӡ�:k�P�L�.Ռ���w����Y�����+yh��Q�f@������&ZUg�ւy��򇠌<UϨ0�j�8�������I%��xȔ��dx�#�x�4�1�[��F /�5cǮĮ2�D�����?PLԶ�猪�C���#�	�34�b�Z�F.K1>N�a'Ў0j,�]�B�5�3��T��0D���:�����A��u��M͊�0�6�Vf�;���ea�"�.B;{$=�Siͧ�qߛ�z7���o��W�i�b؏�y�����E�>A���H!)Z׺�ǭ�e�'���l�hwH,I�Z�?�q2�+<y\�g5�_��x��T
�ڂ�|#��6���L�e��ۤp�G�i Ʊd�%L�����6n,W���E����Fq0�z�cOd2;�s
�G��Wo��H^�W��k�>T����ʫK�uۿ�X5߷��,�}���j�axD�L#�Ӄ5Ѥ炣��?�����}�s�k�`�z{�hט�$�i��I��ݛn� ��^���/��é%�nl�a���c�������bbG/��cl�J���S�y�1,o� q�����lJg?A��1���?:���f���p_~	m�4�$�iX�c'4�h�	ۅ�����I�i�U��3S�������������#��5~�`�t�~R�Ҫ�F�<G���v�JAX��R"����"�5���F)*oVi���82l�D�xr���q'[���i?��<�)�M�B��co��FC@�Ll&5��Z�3ў�:��a(��-�>��$ʆ�r����rU�A׮f�g�%�mͿ���_ֱT6�o�C�'M��?���hg�:��C&\~W%8M���y��vQ��Y�
�B����z���|����9<���D��D�R�L���*�I���Xy�������+����*~���3|~�S����'#���IýO�	�јk�����sֽ��m_IO��`d�L���o�ǣ�D�@]�%�`�A!�L�K'�@�Wш9����ɳ=�Z-q>W���D�Z9�Z�5��s=2%k�:IP]k�)�B��	�UD�e���z��.�EuR��l]
4�Rg�Y��n�����̹#ב ���.\���J*�+ ���g��x��z�y�%�6_�)4$U���]�����
J�8���N�Z��ǹ0���L�W�Q���Q;�e��=���2dQ퓉��R�G��SMY�s��m���cd�9q܌oᵟ_�[p��*����:%y/Z��*FN9��Wt>wQշ��������<�m��N�B�v�s�(Qx��
��V谓$w`��G�$�:(��-l�.'���@��� �,Nr���S��r����(����닙0���K���	�����n��='m�]�늼:���!��Y��ao�Z�7uߡ��Q���6�׽RA;ڀ��Hx�'���$�P��Z4��I��厇�Vs�/a�p_nT|�C�+E��@)��И#c{�d�&?��k��H_),ӵ/<�F��-|�W�<b���M�Oa���FU��>�B�Ȳ�A��P�-SuCr��!�v��K��Ը� �eq}{����H��v�?{�qD\;B>�t7���H�!�z�A)�y� _H?oz+$x1���������z$_�#���l��D�w�5Pg��5��Y0��+ t����K6}�����)r,��o�3v���k~�@��ٸm�Jb%˷8�ee�4�Y�kx��u�۟.47|��{�ܜ6?�o����� \�3񒻾FYԮ�t��H<;B��A �N9�s��������D�5���@ṟC01�0�f�/
D�h�*[$�u���S�ߌ䵜���5��!�S��Oӆ��y#sN�yн%������z���W�g����f<�J��w��|3�o�����F��-;��`K!�B�Vg���	���`L�kK!j���$LP��|���)ä*7�H�g5Ƀ����pZ\lK=�{���+t�t�O+l����iw��e�@�+���s�~]���U��6PZmB
Ԛ7x9�K�5����������ҡ���<C��`�0���t�x2��$�o^g~����NJ��ɸGƭ$�~�٦�L�0P�5!h	!ĸ��oގ���R����k��*s܃u��P)���(ʽ%�A�7���b!�p��Y�B���C��[��9} P�o@�����(0t�K�����7�	�j
�L	��QГP���,���韂P�z�y�v�"h��o��WG��J������v����g���a~&�A���3�>��k9v6dD?p�.N����+wO	7�8y8���8��^�}� �%l�%����!��}lM����lËXp�?&�Ʃxb���e�R����Ԛ�6!�θq��^�5-��M��}Ǝ�(�b������@�p�-����zC/�0pF��U�q8"�a�"CR?��������ߡ�3_�63��t�k���q��rfϊԪd��Q��Qv�I�W
:4{���v��
���c�ؤb(��9:1���&�j���ly��BKz�|�f���dJ+���Ȭ>�%1Z�����7m���g/e���|��^���j�)P8^*&��g��y=�'T9���篎�@�Q��-%N��8�B��=sZ\G��,X[�fYsdŪ�U4�~9����7f�"mA�bX��K ��n"����@4�v���^�=���
��+P"�ײ!_��T׽Q�Y^d8�ǉ����V��M�����N�����3-����,샭	�$�&j�F|)"�i�~2�����Yd��GW{#���F�	�#l���,-lLTt�W��5����a�;~����ˁ�ȱ��	cղ���V֊�	�,M,PՒ1������{]n&N�����U�V�/�"h�?���!�=�N��������/P��V���+q
Y�#ݕ�˪���$��h��ň�琪q	¥<�����]9Q]�,g��̰�]Џ�Wc(Q��Յ"��E�0�-�K��bia����1�j3b�5ҐQ�[_  ��<gmΥud�&?t�އJA
��d;��O�bM��:Mjp��ik�
W,8��0�>�Ǒ/i{%�U��$�E�-�S��U�w@�&}=��00͔V�[O���
}�	]����Y<}]S�X^F�I�5|������?S=�JX�{�Q���U�L��.u�&j����Eo8�^R��$Eiu�}eZ0��{1��\�!��� ����jx��T}>�+ر�h�H�W��,��~T�����6R'�Pt�-��p`�t)��}�ϼY)**���:�����9�U\F"J����C߾(0S**���G��h��8�O���������x���V���]�ǲi��zEz����
�-�o�A�
�!���#��-S�Q�u��&�Qy�oJ�e�j�%�§w
s�߿��n�_�H�	^�~�D��CO�J�^��@����С�꾨ݤ�wݤ���ڕ����F���W�ьi,�~7�䊎
 ��w�d�dz@����S�%���I�V�d���ϕ�.��
UK3�Ӻ4�LS���Ѣ����A��Q2�		]+��7��m~áb���w���f$�R_�퀧qtJPΞF�[�V���W�uD��P��,��s���Y}uH�J=b��5u��Ϲhf�7�1�=�mE8e�-:`���������S��>I���#�Y���c����|��H�΂-����^�{��Np(�oso�!R��'�/Λ��i���̇�rU�p�����6\q�kOH�=�an��~�����ВuwZ%��/�=��5§�~�/J[A�x��.�b�k��/�ʎ�<36�f���H9JhW�g�̥��W�o���w�k�?���dƝL�z;�o�2P��
�����	6��$zHx¨c���lJ.&"m��XmL��s���ثWiV���O���!�ݴg$���c}ڟd��n�Љ�E▝6Z�:�	˛z���2"�V{�i��U$p�b�}(��W��I�7�+]�Nz�#����|̏���6jQG�ܪ�~�]R���+����N�>$��C������>�$Zjvd�jeb����BI9���S�P$���(~�kf�_�J7Eó5��b��%.N)̆ҥ����Pq��	:B�q��Q�Ϫ���V[ ��ڢŠ-���i�A�7t�3�a��F'��� 9�"�A����y#}����`���&�c1�xx)��r�ί�E���}Z����nr�&����`3���G,j6I�kɰP%VzԠ�hJ�3�?b����A�U�m�˷�q*�
"x&�l�b��V.p��3N������{4��!y����i�� �nTm��;)z�b(����}�kܔ���^Z�4��X�����ų�D�Ea~���)���ݴ�y��[�Ͱ\"ǈ�Ջz��@5�����Xс㖼�~S�Z9i��HY�u�Y�"��wg'{�'�8L��C�_�O�9���xN'f�H�5Cbz�A
�n"7����~2�+�`h� lI�}f7� �ܼ(W6���/�):�6��q���@u޾��DIk����s|��A�'��U����XP'��Wp�J��^��/�ʞ)Ѥy�����#ukK�ccM��� ~��p|ܨ%�hы�A���z,����Xt-��\��I���?q=��=!uO�c�"��IݽD���ǧ������+M��BU�c�	�E�����$�pĽ��|xOuQя��@d���0m�>����;پ�/�D�ET��w���?&諲d���%�x=�>�Lx[�k�U
K�Qg����UT�3��iQ��f}���Av\@��`O~υ}�3����t�Ǝ��4^y���a��R�&�)K,_�|���hfk��GYEh>L���*��P�S�n?�?y�X@�g��w��Tx��0T��e��[���8�b�l�(`�����^<A�qj�0Ǻo*F��e���n
�r�B+��q롺�=�zm\/8�%X���L�ܷ��=8����8�7�wɭ/��S��=>��E����Sw�sl�Yxۈ\_���lY]X���A����C��9�b\{2 l��.IޫD_,T#�=����)�k��8�l/���U�f���mXT�n�Ņ�@��3m��v�y�}~�.;�^���~C�b�ea�azD�E��Yt��A���-�x�N�1���W LBɗ�����vW��F�cR�rY�dn��A�`�sV/3J��@lNp,�cVЯ	Qr���F�����:>ѳ����
����(w&Ѳ2#-2,I"��y�אR�|Q�l�* �\5{\�5��@���7����|	��Rz�1r�}��L�����o��E�� ���6�4>?(��*Dz\��"M�	�i= (UWD��:̣s�-��|}-����7�%�F�.�O���;���e<["L<	E�ۋ�� �d��x[VV	}=m �~L_���)W��:���G�Ҵ?FM�J��Դ��Aʼ��]ݴB(�{x�����z��t_�cg�{p���,b�1�G�B��J]�r�417u_V�H����P�op�F�� ��I�P��KG��E����D�Sl�yNN�t�.���<�~�D�"l� =����.Z�ގ�E�8Δ1�O���Ҥ���2%f��T��į�g��k�3|�2�L�h�TF�t!�<��gHw�X���] �(�F~9�b�@���y���p|K���q(x����T��i��Gі��)!��\��J`ۏMk]�4CN��{	z��^	�x���) ?�Xm�8Q=�3N.�(jn�S����Kbԧ�Z�t�:��Cm�V���#g;�6��n���>���l����u�WکT|?�d+�J��D�/?$n"����^��NnL�����|�����{J!�Ƣ���<�^PdcKZn��	w��a&�g����d$�t{]��à��.��y-�mV8�g�ǵ(�!�4�9E-P߇���JJWNVɘ��Յ�U�I�
���e��S�����T�L@���=��A$:ά��P�I��С��O�X�GgnD���$�l
%g��Mߺ���7��� ��h
0y���?p�8�#����\􍺽����K ��&�x�P<�]��w}��d�V$���]a�0�-o@��sQl͐�u�[_��7�2���-fM6<Vq���mZ��;,^"6-<��b�@A��y�����z$�1; ����**����W"�>J����`���B���b���T�6*�=�c�d��:ݚr�a���7�{�|��r�P [ƽ�*�"����J�� �B�1��sP�[O�0����%��P!�g$�^�gG��C����������~�c�{Y�����
_���6�U�F"E���'s(b��9�����d� D��S@�J!?���#Kf�c�ab���=RV0�$*f���z�5uZ��]���iWZ�z?)����ߕ�ᚢ��w�;=p���j�5m6�mτLc���Y+:���FBA���:�V�˟
�7���
;��w���2����� �.��΋ФM2ve�}ضuX�d�G�8�Ж���̨H^�L_|��T��*��������u�.;�0�H>H��w��M7n�?���A�i%����bʍ٥XW@�	'�ë����B`O�*��m����78`?Hs����ɞZ��5S�	#`ix���tϳ�G�Ϣ�,x>bY�-D��E��3�-5ةR��+�U"���/�[�p��ο��a�Z�Ğh��p��2	a\c"��� ��]����X^�md�Ph�۟l7�+��7?δ�&���ʭ��LC�2XG��X� �?���K�RDʛ�\ѷ���}7�vD�c;��E`p4;���@(�{ ��SO�^&anF���N���
q�2���!���J.|�?Ш�E�*I�󃫫&��Ƹ�,ν�̌-�� j�o�TҤ��19-�]�}\L�K�`�Q��6�6��N܇�u8����q�Lj���凊�c�gD{`�h�h���(��^�ֺ%�P�%��u��%�ض�@�����0�,��8{�~O3�7~�D�����?:�/��;foULv��:�0R��c��}�.B���L���O��L;����E�!wm��Kv���J��BR�D.TVz"}�\���g�Rǘ(�00R��?���m�yʉUK�`��*�u�NO�pA;y0|�<#nǗO2r�lwꡞ�.�G�[�
���"���Kcm��t(6��۬Kx��YG�s�ϳ&�H���E~���%"�z���̋���D��o����I�d�d8qF�b>��f��y�����5d8O�"����x'�^b2�P���3�sF��w��$�_����m�h(b��V)R�+sI,^��*�H��}3k�o'�9נ�!P/o�ۤ�]n��2�2��� d�	��5*���u�~k�0�����4?��$lZ��d���Z��l�v��0 �0��V�_�Ԍ�������}��:/�����=B�夫��JD�(i�b}�SC�Y@+�������.J2��@Y�C�N?	H�m�&��)]6��� ԪK�(�!��lm�"ݙ��\����O�o���Q\�6鸉ּu�0ෛ����0%��دڞ�F�hR�}�G%�/g�ִu�E��G>��X��Mqf����5��ҋMJ����MD_A��;$Bj_��Y-����-j_}_���*��	��?@Q5�UhQ�~c-ev��:ׁ�r$(��˷ރ�xs11:�=ͪM�E4����[�������%}��g���ρ����Ցq����T�h����^P��0�$���gXB-�&�.�8��ܥ�}�C�·�&����a�w��'�����W�?H��U�k��u<�����A������Ջ��p��C�G�5y�~�a���H��D����C�˪Խ{�s�e_�{��yx�۸{�hv�㶨�p���´IX�'53c��yã�TD�q�� ��e�ż0w����FI<o{�0�eAg ���#X�[���5!��U4u���}�R����f��:e�Pqw"�;�E�2W�X!���I`�U��sZ��6�P�%��Ũ�۪&����_:ZJ���-�׬U�nFhT�O
�e�lN��\�Ts-�k�'�12|/� �����=�Ǹ�����4��E:`F�;q�N�.DS�M�  ,Fj���k�-(��a�1�|�g	�"ACQ]B�[pc^+�k�	��pk�!�L�\`g�O5e(����A;���QV�>B�����]�J��i���R���GaO��qs����b������f��	=����ԣ45,D� "ι����J	���f.�@$�*h��Ņ)	A�ϸ�@�����3-4��>�sr1�v���SKa-<�w���e�yq�0���+�-�[�]s�}�d���xsm�Xev�1���A�ۈ��-I��A�d:F�7w���"t:�}�L�� F��-�$Y��"�Q��M�n���-.K���qzXޝ>��@A>J����m�P����D�����E�tMg��ů�c)H;�R���sD���s��0�0�fhdU�u����G�/ �F+ȜbYT���a��Y\�6���f&:"�nW��x�/��[zz64���T�@��z����A�z��m�`���-�F������+����$�M­	���هu��|ʥ�U�y_B�+$I3yT�����s�_/�ܿk�����zB�18�ЦF��M�f'�K����\�~8�ќ���6����*��ʘ����3�r2�A�XRD%��y�8�WW��G�*�k���l5��&%E�Ě����&I����cMb4�h/�&����J����w!�K��C	f�L�ťa���;��8
�eĪ{͉����T�)/��s.Xe�\%+�@k4|��~4���c��z�
� 4S3�����]Ws���T.��&h;�՛��E��]2a��SI=���ro�G�6ch�V(�0:s:��D{^���c���T�g}9<B�1($��}���Ω�y�D�H} C��7{u�@o \+\�x%��cqK}F�ņ�,����ܫ�y��s�u>�GyK�v�H�vv��|�"]�3vDif�b�ުo��W�kUܽ��$��w�!��';P�6��A���Z���1+]Ώ7�t>�&�������7�B�'�y��6Ѐv�/��nP\Tl}��t�܊���Ǿ��,4��S�9��DĎ���f��r�0Ov+����.�L$��g[�W����H�\t����1��"�DN�f�����5���>g�!ΖZͩ�o�Y����P��=�3�6�i~e��_6�S�[BӋ�7���U�d�c;�)�뽎�kG�>��_�M�`���a�U\�n� �XMG�4Ɉ�C;+W�����mf6$����Yh�Z���#N7���n��=l�I���C�b�'8�_)�e��"¢̹^�՟$�O�X�� ���1������+1o`�G/+��%�";_�w�>�����)Q��p�%�a���ST����G�����mˮ�X�@s��~���z�f=���8PJ��#�����(-����`H�i�����v��2�<6W��*Z$VT����ؑX����J��;˙/y!����Q�FyJ�D�c�~��o��se�ա��?����Y��Q	�Q�?���g�������'\��P'A�n�1	Dڶ�n���am����xc���Q*�Gn��k'�^�2���T�=g'��GX���Q#h;mv�F.EV%�~`T}��
�
>�T��k�� YWe��0�AKMyٸ��Mݣq�%�e�¤��w|<�Z��eI{��a��l�EOc2��*D>'O�~���ޯQ���j|v[���RpH�J���"����ߌ���.��q�>]�#�2 RQ�.�������t��Vkm\.W��2Y�Z�����iD�7*]�;ܛ�'��2ߖ��v�e5�U������L�?���^Y昪���Ln�M�Q�bZe~ӣ���q�,����dD���*���vGU���c	���i�״`��}4��Oi�\;
��Q��f�p�Ǎ=��ӥH��&��=OfGg:j|/�kRۥ�~�#���Ҩja�sJ���ش��p��x�d�+�s�4�C1�!��u+^l�����呞l����ǹM�z ���\{�Qr�D��ÿ�{ݦ�JϰY�����`t�[e�:����j�9��"L�2c+5�#��J���K���F耵�9�H��7Ku�$ �(�a}h�S:��I|���;�f�_�U�S�O��O��<�$5�a�f�~�G0�ֿ/o̤�l�,0�z��{t�p� �!�5�l��Q�#=��@'�gKr��@@�o�aR�TϪ��~��N�-���<zf��4
��Ӥ}������$:l�oЩa�V��yE�m�Ӡ}J�n��x6��Nv�B_���c�`���i�6�w+�n�y���R��x�����*�wPCV���������/����e�@�XH��anq�<j���+��n󖌓�	σ�;͌�S�׸S��T�0�D���K���츸�[�i �"Z����M�����U����*��r|����C-z6�&�|�]�e��x#�7?��mM���Mdt�-}w���������#�/���`��l�&W���l�}r��5�t�]�;J~�gT3�)|�	�~�q��o[N }�H:/��x�83�n�0��l�x�O��kAd	L4���d6�b5/hO�u]����~�����j4HH9��a���0�r/C#�>r��W�X����.�:=�mj����Z#�i�����6!�4�v�ʬ��X�����+����Y�Z���˧y�
����<��V����>䣵<��>a�˗�JXz���5��~M�n�q�;.�?�T��n����Ts�LLR A���lJ��ogKʤ� ~5��~�bj>�D�ߣ�o�od*�2L�i��ͩ�_�z�9�pa� Ӊ�����,��̿H׀y��������N?e��mC�E�#�{-��Q�^þ�������fK����t���lʲ]�ߔ3�^���-d��'z��~|����)[��Ǎ����h��v������������-T%��7��eh.�I�"J	"�N�W͗�4D��jW�H��"�5���J��I��׋��0Q�=ST/AH��M�d�\�$�R7��*t�Gwhi�ľr�bD�S�l�&sP��}ø[�^��\�ωw7�X,�ޫg����Z�q�Q���Ŕѓ�47z�V�_M0�K����p�9�W,O�@�"~����� \;���Y��K5 �2@g)u���ϐ
�Y&Y��+9AP�N�N� �(��-H��"�u� P�ݡPzC'8�4�?`�U~�X�MQ�.�t��G��``�J��w �\~[`lӫp6Þ����^e6F��.KW�M�zg
��V�7�oś�@B��g+�*���^���mߑ��|VãT�S��G=����:�!�2��ċ̛���r�-�JI������ٙ�����Woxχ�,��'�ۍ�	d�9�^&�=Y59�xx�Q:�I\6V��^ٜjAZ���o�:�Dcς�H2K(�1ߧ�1���������=�0�����nQio):;Z��ɪ���E����#Ӗ�f�=�Z���7�W*�X5��AN��Z�j���#�e�����.�/�W�aP@P�`͂��FG0=-*j���\��
h)�iق��㊕T8u�B����A�yRaZ�za����B�@"�+-d�L�7��y%�72\_�"1�3��%��=a���S�[��!�C���_�s`����?�۩jPr��A�
jh��W	(D��s��ِ�/qS$A䧱�������o�2��#��*֛N�L�.$�C�y:s�:K�E&����"�E*&b�ֳ�u�#N�����J/��Q���ń��'��U�]�~gø���M�H�8�Y��%$LAV����2�������l2���e@��>��p�f�i$�2@@���oG����vEe��������OU<����)�C"B��j��ݬ���>�\B�*��!�v�=,���:�i/n�ƈ�I���L]m��	��23��������<�n��Y�ޥ"#��f���^L�r��'RD�}�8r>bV�>�U�2�u6D�:tw�>	/�H�F�t"����A���-�Ƨ�&�i���̾������aX���"�f�>m��z�Q�T�s��[Ш�-LI���>j�׍���[����2mg5��]m�j�'=Q�h��i\�&�������W����?JW�ҡ.���+�оp�����
�quu~w����^�;�l�8ۣ�Yڒl2E~���)բ�k�X���
	��6S��͎	�K-��r�֥VC�\[�\�G.<Spd�4���"H(9?��R�@7s�Q�E>C/c�{��Ѡ�7Y��V�~���yx�k�UI���	܊DPS3��J�5�H��zcU�J�e��ĵ029�w��(�\��8e��/c���]p5̤Y㒄^�^�������BQ�.c�hFI������l{|X�b���.����u)��fqV6֑��r�J���/9.��#| �>n�AG¾����L<�.�5�	�m��p�@��m�U��pyY븲��t�7;\����$w&��v0Kl�=�
zR6@�^���Ȩ�u�V8�9$!�N=(�ߋE�*H�r�w��\��������΀W�����ۇN�������� K��������g��ǻ[��Ç����}��T�u��qRY��r�����|��Da`vcf�r��l��Ov�j�M����J�#�S�c+":���F]M�jt��$��@�^�]d)L��dh�@q�>���tB��Ӗ�* 4&D�:u`�����>��n��� �޳CKЮ�ջ��!��`T���8Ƭ)�A�JxGO��V�K8���%�>
���]���e�AK�1K�X�1f�^Y��m�2��3�v��>���D�ם�?m)��wz��o�v�(�������7&��R�^
��A'���)b�g���
���:f ���0�\��c�	Їg�aX���l�:l�ؚ"�����V��P;1;�=�u�w!E�w
�qT�`��r Q��WXc�����ד}	\:"s�;z5Sb�8�Cp.6�6�L��Y�K�U(���|���(ǳb�6	�s�	��@?���}�����ͺ��Jj,�9/�]�]a��)�tEkVHF��>L��u�(��~�	�6hAB��~�y� 0��+$s�h~>�I���k$�����
�!y%5�.�gN�#��"2ɉ��'����_=77�C���������-$��m�\��VZ7d�$�y����J���w�����s��97Y��'��]���f������D��G��t�F;_��^�����=~�ʵ- �F`��|�x�x�a�C�
j�D|���=3�"��m���T��ZB�X\�&����4�QIQ���A��!"{����JS4����Yy?/�g��f<0JR���ջ&�%0�d�VΞ-�0]�d���-ǀ?̙�O�[!�E!~��J���W<̡�E���,R�9��'���TM���}����zvsæl4�^��Q�B�2�^AU�$��D�:�K�{�Na�
te��f� ��5��w��nmK�i߱�5l�ӕ��8TbO���<�
iQ�G��C���F ��u��U��4_NCf?���`�8�=�4'�jx}��z�!@�'t\_3��^ߵ'A����er(�,�Ŝ�|�/Z۲&�xy�m.Qz-l\^>,:6���<�`�"6������`�+�%�-��s�۾��ҷ4�:5�"M�%� �T��-Z���0H� �rء0���?�t
?�2�5�_�/�n�+�e�{��ʺ�p<ߡ�7O�5�c)��'�m�H
8��ʙ�<pY͔�A��q�5;�F�3�iW�֭���0R�,���apb����Zf��,ؔ�\��w�� H5B�P��;'�Ri���s~M����z%t����.�r6g$L�&�&E*�[��e��V��&G�����~^_$��*@���/�LӚ��Sԅ�F �IF�)����]y��]��~�}=�M���(��Ōf�3�iy:�O(Uׁ�hԕo��h�! |��a�h��[1���,4rPL�g��s̡�:eTV��S����f��^�8��R9x"����Ř9	�	mb�����Uj:��{gH��jﳋ۴������ݫ��
�ʲ}�/`��u� =t���(��M�ZY87��¢{�T C�� �L�������2z��q���4;p��z>.�eRim�l$1��v��o�o��_Ÿ����#x	U��ԛ��F^�K���wC���g]�J9�(�������Ī��)���tҖf���@��H��43��^�V�[=�zT`a��։$�[��%�~�u0&�e��֐JZ&�@��^�[J�����Τ<��N��4˄s�Q�,a.ϰ.
��������tb��Q�r!��/���JCj^� ui:o=��r�<�"�u2S�֞��#n�G-*����$N��+�*|1���*��t�o���s�Rf<X��}����0����H_�DZ2b��*3��n��	6�{�>DK�}�*T��qNmy�L�-�-���h;��gR@��6}-ɃB��:�==m��#�<��Y2ν)���gx�R��#�i���z������˄<�QXя�a��*��n
��$^:xO��o�hQ{�YUrْO�u��ę}�a7����@��3(wc���q��#�b�݅u����dw_�&hǀ�a����k*{a�v���SV��y�O0!��k�]?�k0��!G�'Ŕm�����֨.zaĤ:ㇸ@��W+],t��=3�*�g�2��_��cg��z�m�n�+�� ���h�=#]8j,�S��2�A͊���(ӱ�F!���}��[�-Z��]�G�FO��پ���I��7a��ӶOt� ܵ�HErJm���21��y5(
���f	Gvt���_g����Mv��Һ3�,��)�ޥ�9WrԦך��LI'� �� ��Rú)�+^2��}�p��#�Ғ ��G�9��/�����܇o�/'� χ��Ck������}/L"Ϊa��'�!�a[�*�����km6����ΦA.�\@汰N��Rp��g,um�����1 �5V��!�ۚ��,7��4�l��XE(^�,��]Όy�����c�q9`�*���U̍ŋ� �-�!�˰h.��pi)���使��+�� K5hhSRaer��I6��54��p" ]��^�	R�����۩�r|�Vz L~?όv��VP�6� w>�]�.l�3�R�j��ԵoXGx:*_�*�wM������ D�K��� ��$�|��s�64�DP�Xk�3�i�M\m�F^O_Co�_��|�'chy�����6T	���Ȥ6�k��3�4�����g�Am v/d0z}�{i���^r�;�w���������� ��ϝ�J�ϓ��g�.C %�9��)�C:�՝T���;��S�\�Ҍ��)�J��7�t#q黽ۮ�**+���삩�|�bx�[�g}^�����ġ0*����f��7�;��C���@-��J/ݎZA�����y>ʔ���-���ʸ���mA᳀��sR����$�|6�4;K_POI����=&��x�P(pH9�:
���]>1��km�V'1�w�G���Q �p;�R�S��I}�{�>�aU����
�\k;L8��tK�����,�{���I�~,i� 7�̗yפ��P�
I��� '���B��3:���M�0	����ٙ��&�:8	�c��:7	��a��_������M���bJ���<x7�������Ƚ�iO}�(o�	�^ɱ/BRES,	%7���z���8^��l�4[Ǧ�oN��H�2�	`�ߦ��.���¨�8���W��m�:&߹�5�o��z>�����2_~X�6��c��ΖG��>��3���5��b�e�i��/�C#���;�=f����^8wQPה��p��n���o��	�9��nU]�S�(c,�v�]�H�S��2}Ɠ�7ģ�#(]��uf*��J8���%�y �!lq��~6��m�pt�-��(uZ�@b �9�����	?ao�.�wo�P<�w¤	T������{��`J�OW���2O��P�.��܃~�!	��D4�ar%�0�B�K}���rAH��� I˲�^�>u����i6�9�������N�m�T�ۍ��I㽑g�j���SOhd�\�W�c���&k7���ZK�!ng���v��v*�	U�T���B��!�n�w3P|���S:-"D��T��̚���	��}l��1&�0������J��F��	�}�ܴ��rU�[�E*�
��� /��5�~�3��nZ�i����&�4��h
�5v�\ܨ�)g�PH�*���d��4�"���$M���h��ON�Rm8��KC�L��p�BP"F^qJ5��4f<�&viI:� �B�]����R��Tn�ٓ�� ;5b�=��}�םQ�q>y���2T�����r�RK�7����d���/�"���EUD�п"m���i�|�u�tn��S����.F�4�GOŕ��ux\����A�m�;gUB&tyv]�Ҫ��\��^`X����y��(��RgT���J���ޠ���w���e�ZMC*�����s�ҧ�?)U���Q�q�K�mx�g��G�����t'���(�uA��l띤rp���`�4����Ύvh.s^�B��Q�J�%���qS�d�i�遵�5����i�F�8�Nl�iՅm���^�]8����Łi壂'�IG2�s>u�e�.^4�s�e��}���t�[D'v��/ؐE�;_vｒ{��c\讄V����U�������d���pЦ�����ݬ����b}Q��,$�GU*euυ���������L:������ř�l=��Ȇ�6�w�^`��ѥ�}xz}���i΂p���I�d����e��Z��J�EWV࿔�ǅ�hQ�Jo�@���e�2.��+6G�R�����B}�F��]w�$�&������fŶHH�iǤ��mM�*�� �$��~�m��!��iE{�H��cW����]���h����N�Q����^P�I�-d=cz�q��p��:�|��j�ɠ�YNj[qU6p9�06��7�d�P��N����j����k������9S*;UT��WG^�~h��P�p]�h(�bܚt1�.}�K�Q%+���8���G�g��ִT(Cc7nJ]A\*��[��z����w���4nɬ��$��\����&XbǙ�`�0%���pb�^nju�l�ό��e�J�����z1�ͮ��G��>zS���EQ ���*���	"4�7��r�OKP��[�)�V�9��:|�� �ԕL��C�S�@Yoьp>�]��&ZںT��b�z�]McZ�, ���?�2腯�b
�	#|����Pߜ�����l�!�U��|�)��:���m�t��f:����� ���U{��*aU�E9��P���.GGC��=5�u����S>��e�ug��45�5 �>��	��fP��
}:֞qa��08V-���^������iC1vq8�|M0=_6�
X�:b]3�dS<��k!�!�MH�(�	��d,���@�<��j���4���G_x��,$�}z��G^�s	��TH��ي������S��w�F����MXωk9f�{�q�R!Q�\||: �f̵p3�C�ѕ��D.G�^��k�w��mP�<���U+�c2`��Z����u�نW�:O���aw��#/��i{�st��PO��,()�2l������.���z�	���`��(�L�^,^��xz�A1�����K�^����`����1�
}f��1PT�	������(��(�����i1 w�� �z+i<-v��5���}Q�H��m��gH�!$c�y""�W��bt�toQv�w�p��rttX��'���
O�ڭ��J�����|�QRk��G��Y����~����ޭ:�+�
g�����E	`�s	�ȝO��k�v�f��8�WN_��v�o8��Y_L��"�>�W�$���S��h��o%hd$^�VO#HL_Wa��.���|�+iB���H��1�F���_O��A�'*W�٘YQ�E�Z��QM��b�m{ ��7�Xr
�ؾrU��3��r5�ܓz��	�~Ib�(����M ��'*y��r��U�K�|j;c7�'��ݚ��K��D��#��9Z9�x�X�ܗ'*��#�)�>`�!��<�� *�5��a�夿Ь��L�Q����*���ؔW�� =�i�Q��D�w�+��xD!��P&_6k��Dz�.V�$ǚV��N����eY#v#�A�YA�Tӎ�Qu�!�I:�>�h����l@dV̽bd����}����j_��Ƕ7Jcm����)LUu��C��o��,�����h�6Z�Q<��R{�IA��ݘW �Ɖ+Xn���(}@��E6�̑<��|����H_���<bkt��s}�in[�QNFڐ��c�Ϋ�b
�Ÿ�!�����U��X�=J> nYl���("�J�ɾ���==T���M�c�Si�i iA��5j�i�r��,�T�K�lx���-��
���7���uL��wg��0PaoN�KsA0��2!s���$f2�u�����o����E���szH:_��ڮ�f�i�,$�(�[��x��& )����U�
�v�k�k�E�P<�'��*Β?z"׊mΆ�?em�?2�m�*���> bD���g�/�-l�N��<�q��δ�2p"��KA��p�Sۑ����~�D�P8;W��K��r��r!t"]!�E;�*�Bj��s8�r�������/�L-)-ҧ��Ɂ|0K��㥯7��3����2��*M�<ݙ��F��s�=��#�$/�y#�B��HI�E�x�54�Hc�)�M+z]&��X�*	���V��HW��۶��ض������%��#c-���|�Cr`:�м�,8���~;�w�8�8��>
Kz}צ1$���h�ئ�s�	6�8����y4��A�O1�������1�aod������A�O���G�S�j�Y.����}{ާ<�'��n�S�j:��.FZ����=���M���g苿d�L�_Es�;�G��P�Ghg���}��2j���(u��FP%K0��1�4��ŦhQ��l���(A�=����>�g��50�bv��=��Co9�2|ԥs�Bp���7=đd��;�6����Ja0d�dP�b1��(�T��u���
}Ny�[a�2'�:]��D��� ��*,��r|	:�)�<��L<L=lZ�����p�Z�h�Z5ѕ	�ZVR7ۿ�e��! ��*ͮ��5� ��JDj	��Y5�H@�0���"�ߺ��0��N�q]/����i�F�����:O�X#O���M.z[�8o9u|x�*�J3:3��4P���a��J���)}ϣ�IV/���RU�Py��U�9pw����I����͇��p&�N6�g��:���&`,��
�W�11�鍶6�1�uňS���#�D�3�Fg�h�{��D�R{�%߾:H��ǃ/t�)Qv^>Mr����js���K���C��K�9�(��	�?Z�[,k#�����=�w��T����/�O�k'����5#*fa�>+�i�%��5L�J��O�W� ��"-~ϫ[�Wc^�伄Bo��=3�h'�<�_l��G�C&�b<k�BrK�>���:M��XԆ�_\���a����aY� tV*N���[�)����&СL�\�ړ���d��-�f�܁J#E����l���Ϛ��J��&X���ǃ8s��RÇJst�fBc�졊8#�*�G�k�I�q�4>��"4e״z=�R����d,|�>z� _���V_⹽�~$�Ul�rk�E=,US�,����S��1�%��Ԑ��ԩl�� kCxk~b��F��v��Bݭ:n��CFO0,�����XܣZV#���J(��	����_�3�ٻ�
�X��S5�!�V�;��1b�S
���QF�: Rʄm���2)�a�vr��}��ܣ�O{	�Ce�p���c��Z�ۜF�Gx�3���Y�"%dn4�q�����Q��$M�D��J��'������%��f��j���1�a�o���a�N?`<A� ���(a����D��4S���؍�&@����{l�j�8:�Ŝ������y��o�=��;v�p����M�M:+		
�B�o�V�t<L�9ư(\ڀ�tPF�A~��>����"��ߺ[�#�����MƂ�m�-�ήb��aa5�[��`����f9��v��L�B��Y����7\�5��j�:2�6�,MF%L�C����`
�<���u��/������);����
� V��b�wX� �6�j�����\�Ӕ���0��^���RtO�^���N|�5�h��L+>���9��@|���1���A����uJ�f��['����A̅��G�!�m�`e���E�ip�J���kP>�y]�6r4�*$��g�?�9�4�n�t�b�d.?;�'��#�}{�4���Hj���;�zB`������\_��hLjH��Em���Ptc
� ?�N��'G��� !�<���$�ǐ�w�7}&�.�ep[�ؗ�����n7hN6����������XKGV��C�*D��cU�+�.l��gORݧ�T�Z�� ͹#Cf��>�8Bԛ�aE��Ʈ�i�T��z�� ��^����`uZ�	#�Qq��⁌v]���~�x}�I�8�I���G�s��d��u#���s���"�T�%��q�V�mx-?rބs��1 QXɭ�J1�c<�~����Mf1��˦'sf9�ú1*x�׼�����8LI���:a�;<�\K �8��zm��Ja�51'.�AH�7�z�e�� �	pBP�P���]��^�Rn	���M�P��^����-3C�c�L:�c�}>���.�8�b�'��b#��@;j��,M�����-xM���F�awӂ��Rn���ԥ���S�B�t�	�Њa����z�̷Qږ�J���~l���e�x��Ħ'���~��|�Q�z���c&�M��n��+5܋�*!ИƮ{�����Į��s�yY�)��˻]E�!=bB�����A���c�� !�^�P�"G��O����G�L��<�'0Y��M���噖^%cL�f�)�w��-���;��b�ү��Z���%K5�Adt����y�l�5�>8Y(��f,V�q9y�"�y�B@e��5�~���L+�h��q��Id���D��M��o�E�֚�ƀfQ.��/�v�k�]��z��(1�8�.����Gb�,���Y����qB�$�+�UZJI� K�5��R�����/ݠ5�~Ϗg�0�T�k�����!���Cs��D����i78R����ۭ:C9) ���v]r�t+jV��1՘(��aJ��j�Z�� �60���bAy�{��h8���D`�g�Ƽ�>rr��ʴ��P0�i���T�&t|>BV�kD{�o��B�h�J�[���$8x*����|1a(�Aj%󱼲*�M����?���tdS�Rc%�k�t��x�h�����������~#�u����M߂+xl�H�:�q����hy���T1t����W��@� �a��[��t `"[BI����t�e��U��-9i]�sNX�U]��#�3}>��c�֪:Ta"��H��Ϸc�4��J�串��h��̌����c���c�ծ�r���Z�3O�ɭdM.�W�e�J�Y�������6�|M���Y]*�;$���8T��v�M���#j�}Y��]\��D���CvS3M�T���@����y��ډ��InQ�D��r���%D�<q�H�5VTP_�Oݙ.��/�\%�{��G'����\+�Xם���-��Qb�o!�^ѯ�TP���m�P;c��������y��\�0VTP��	��� ����\n)+�O��ꈹ�I�#Lɸa}Ň�9����#�kQ���*x�
�|.j��fX����{y��&g�a�I�0�k��J�Zl�]t�'��(��Xa��w]LmL��3�(��Ó��H�~����-S����^�r�����x���5�QT��'aӗ�d⿷�l=��"�K2�L��Iv���yDz�>~b71�QXB]�V���!<���_���~�iJ�t����Ͱ���Y�G�~�*����W���yL�!�2V�W�@4=c�� ��;Q5���&��E����7�4 h��E	&���k���N�99(%G�������;z!
�7V5�)!œ҄�����̤$���P�X��s��/�>8ܲ��{K��T%���̕^*_
���"��摧P��CEش�9����w�^��Ƿ�5�8g�D��}���1U��/�@�d�3B��z֫�Pa�x|O��b�vE#���:TŹW�nĀ�B�x�{�@��3s�נ;��oE<���!��\�Q(ɇ�q�m�A?��s���B����nR�f�kY����:ٝĐ��XQ���Do�x ��D���?l[>̈́���i��.�A��I߼Y��u���&��䩮�8����^O��c�;���!6`����I� mr�b����9�f�̯�o� ,Obĺ,�>z�U��v��a˾݆ ��fă'j*���t��n���͠N[L��%T�"YN���i���BP�^{ %Ǽ�(�@��ݑi�-G�Q�|���5(�s�JL�Zx"nPA��s��	��~��,n�������uxZҎb����+r�[Fh}=�2�K'"�0K��DT�[O}�1�n�O:�A!o[�=H�&vk�@��y�ן�=�*hxz� W�%P����{��]H�+���6R��$���Nu"�-�fR{lc��>�r�R�#�_-�=�#�Ǻz҂=�\�~K7�m7���}>X[��]��&�@Y����TM�>� (i�|$i͏,Wx���Y�ؙ@��'6�S�f��ψ��p��7��C&2^9�a �oʞ�8e�d� ET�A?��3�]L0�O!D_�މn�'7�˃�@��]ԩ��u�&[��:��6�r7>&of�
�@}
m��eޣw����9B8NⲰ���ގ���6
�\[Q�B�r]�O#5�W�1r�{n�����0����k��i4� ����Ͳ7}E����I/��:@]����L�.����ϝP�҉��G2�#�����7f��i	���|{�j��ܥ�����E�;�Mo�qr~u��*Kr�(!�t����g����=X\��1ޒ/cu��j�������}�:��aW��
c���`d J��'��� C�To	M� �-]/������<~u�W=�����Z)���w���O�R�x�lY�yu4WM:��Y�O�T��E�w,;$<�zT"�E?�I��H����-#�| �y�s>�:��z�k�|�%����5
w}�m�`���:����]y����Җ� ���f�D�m� 8*��X��.
ᔔL�r5\��w�;߹�b+3�,c��S�ÿ�-���_g>��wk�~��?�0�A4��	��p6���<�6� ��o�w�Sn�M�
R0�n����OS�k]�Ƥ2a�v���p��N��L��ia�L��[�]UG}U���`�Vs�N� k����HnS�!��z�z.��n,�3�	�	Ф\[p�J�9��4�r2�����&)� M2����y�d_��C��B����U�O R���'��IAB.!�Y�c��#�s�?F:�+�.����{�4"�����zfQꜿ��'7,��2[��Jp� �Th�/\�2�tr��<J�Ĩ��4���X��ʯ����ˍ��Nq��?�{�ti�j�o����p�V����a��#�� 9�g[����D���|�I�LK��!�_⾳�i�w���K�4�=]���ށo�x�?��G9�2T�?q�T���"3Ԝ�ޕ���!cv�}���1�=��E����Կ��e��i]f,W,�ӳ��\�����������+��B�f{�9��}>4Z��ݻ��n.+�:SF�� ��;xŲ�n�p��fUg�'��W���W�����t��k�̇X_ �wNu.��Jq��J�$��(D�OŃ�}*IV�=�����]�l���4h�d����a�)I�+��<��v�=d�l�ŭ�眖 �7N�Yes)���7�盞R��R<�%c�0v�C�!﾿P0�Sg��l��>v�=G��C>�%�����]P`_"T���	^k7���rր��t�E�ϊ[�%�wqa�蟃l�7��u�7M2)G��B�!��Zr)�rNu�!D�^��;8Yg��I/�"�B�~�Dyڿ4�9Ĩ�ӷ� »����@��9���.,���|dO͔��������%�9򵓬���R9�`��?p�{�4	�������m�}b��3���8�2 (JD�ڞ9U$K��Έ�b��.�Gl��s�/���R&[��K:J��(cj���̨�~�Tm���`�6`ޣ*�%�����"�.K�ʇr7-�����~ۖ3��_Nֳ�1a_GE4E��O`3x��@U�	�6���V�<��T�	�f%�H܆q_C�z�2B\��%��V
x|V
�
ۣ��c{/[�/��$d��&X&S��":Ի�:I� |�-���>����x��=�C�O��O� �� ���wP��vl���8�pt�c\�R�O�T�&��w���º����jü�{b;b��AB��ұV��1�=7�f��?/�{l��Onr�ؖ�_Q�{<񀈍w]�x}wu!껔�R��N�
��?oP�AI&�+��T��;��Q(�ɹV<~�����n���BrS=�����<�
o�8��H?-a���P��ГŚ�E�j<���$�:���.�S��T�<�(���q�|屽��P6zR�1@FN�(�.�v�������;�d"�	��4��$j�b�
�m�S���=/����M�M)-˶�l�p$e�8@:�0�09BjԽ�PA���#]6�S_[��)�J�e�}�;��K<٩��Ń6�s�y��m��x��)������
^������`�����A����Y$����S�X�6$���*/	�su��FH�A��gvJ��v��cdQ�{_>`�M��6%;���7:�!�S2�$�����.�W��x�8S�ץ��ğ�ޓ:��*}���s�G3ꄩ$H��Aa'$���:	ণ����vفK&�r.��,w�i��PX�1L��4n=�G��ƕ�''��XQ���Ӡ���A�S��D�SN��¹�x|�����5|� B*,�Z�>��r`��d�/��.gc7��2���Ѷn��F��^��� ��S-��@���M�;��t���Vf��V'F���F�v��ȠW���	�2�s�
�PTڣ@�z�Rj>�'�����'��Üx��*���a�q_p�
��L��}y�c��)�;���n#�����0Xj(L��dt��ԙ�a	л@W���0��Y�8%[_���etƹˣ4�����|���kā�m�H�� )ue	���	�A���r�LE�]�j��.���)��<�l��p�J`��:C�����ɦ-௜$�74����>\ﾑ�[=�p��T�i{V�$����i����u��r���(*�P>/��$������pEV�V+5%��U_���hx���н1���΀b���.~�H.`�q �6�����5	� ���'����P{���M��F~�W[PwzV��8XHH^F͵���*�Uv���5-��կ:��D�Y�F)�Vv C�x�s�������N4�u��w&ӉR����o֤M-k�lA��E>���M�y:sY�*��/�Z��~b��&�۷�x&!�-NGr'���w�D�J����޲t���Uy-�"6:6�0�^+,9�;�*����$,�*3�3o�9{�YSI��w7�'s���`#e��J"�Z��C�QEr�ɏ.�����.Ȅ|>��W�w[Q31�u�����-��`$Zg���ki���.�'v�Xd�������yW@T�4*�ڼ���+ x�� �ó/ك����up��<�/����c�����>yW�	P)O�0����i�R%��ċ���9)Za*�rUSS�P�4�rzg�=�o��aZ�005���d篼b>]���^*R�2�nj	I�W2x'd�,�������BLA2�H�S\����0�f{b%Ȏ���T�wy_YN�+��ߚ*sg�5"o�\���uE��L�H#���#C�(WP��VbW�'�\��Li�V�ʩ�:#�J���e��X	ņ��ԣ��g��9�������o	q�IfsZ���-w"T����t)����e�!�4��v[�,�Ն�:G;u���H�̮�@?����}��/ ��;ǉ��B�٨�7�z��GC�U/^�)�'a1�P��4:<�9��R�V[��C\�Q�p��
,D���&�(��,��_	R>�lB,���E����\���D����� fY�)����腣�(����%�@�y�ă��^�}�\�]�	����ߩc�N�U����zᛳ��h��F��	�bq܈��jg�Y��o�
� ��f)���)��N��J�̐\�&
�À����O��8B!�S�[�bS���\
��hU��5��½E����X3h���s
��	O�gM��L��O��Ak���eAtz��ѲE�AH��Oop��m���`KaK�y䱭iwW��E~��i�Ҹ�q0 �S�~���}p�,�*��
��.�>����4t�����Xi������"`�zQ�����qM�ڝMj�^�;4�5BZ�,�:��_�����S�� �񰴐�`;���b� ޜhg\Թ#*���!��e�	���=�F��Q��]!�~�cw������]�H�O�ݶ�r��z���ⵙ�b��~�����^�&�Á�s�яx6$N7P���x�ݝ�b��֜��a����j�(�0X�I�$��?�u]y��i;{��Jy�x��d�4���->�mt� Zj���w���;�g�cz�x���#��Q��F��v��9����3�)�6���� �~˨Bº�=,�C�Өf5��W��A��&�ʆw�6,�m�O���`�5��EP�!�$�1�R�o��7�����3� ���
���p�)w#W�m�	�`�&� ;U���8��]%�����V	����M��^ܗ*��,�ESh�&(��n?�h�^�Iw�;4Q!�͂VGo�h�����ɹS���t��q�w]3�˄��L�6�f����ڌ�U�]��fx��q}���3n�5����ԩ�~�Z�,Ӑ��C��Sh��.�w7�iSV��K @:5��u\�~D�,�R�琈nf:\�?�M��TW�u	F8dgzMc�Ti��P!�)/̋`���X�Z@P�b�2~�#"bF]����OPE��ҾG�Ǭ
��%��E!Ȳ��Q�C���_�Y|ΠȶR���}��|�`�s��|���`��y|V	���o �2e@ݡ�I���-�:}��JCL�}�ؙv�����.T� Č)�ĝf���Q#�lqA��5|�r"���
(��%��"������e�W�j��&�Fpg4~q�S�*�h!<E
Ѝ�~k�X������AB&���u�n�o��_�q����_��������G@�~��-��C	2�G�#����0�������������JC�\Xcj=�a��b�Bw�]3���g�p��~ڑ(�ha�I��-#a�E�py��Y���:5й�����g���B��=%,�G��J
�}��C� ѳ�x!b���<�N�a�8��	P;Rw���Y�U ܶ���0�;M� Se�^>TVy�ѠcV�*!A��E���	B��+�H�/��'8UA�"�ޓ��ܴ?�<n=�-�*�E���M,�����#�>�yJdS�h�-�k69��55�������i
L������y5���,t�;��J��E|=�ۈ��p�O�O��#�Ҷ��j��4L���Ӭl�AZQ��]fT%Y�b��&��۷R�x����CY��\�Vf'V{<��3)�Y�17�e��l���Ĭ��%���lDH�zs��f�$riҙa���EaH��F�<-Ln�7ר�G��Ҿ��L���'\V����Ծ<�&�s:�t�u׎i�]�T��d������]m�k�s����s��?�z��'�vڰ>�'�a7�2�����&�:��
Mf������y����dT!��Pq�g_��&�!�{^����h��������i�Ѳ�ʺM�vEx#�r�Ǌ�R�X�ۊ�]��lkv+\:i�Z�xӜ��}Q۴�ٽ�3�1�OPԫG��.�)�*K%>Y�#FI�()�TWX�Z�u*Q?�r!}��J�_�U,��\�>�+�Vǋ�\�?��eC����[�&Ơ��З�z�X�.��|���,��,[�OTJ��r�*����Ǜ�zҖ��ߵ�Q���-��"}�1p����6B���@,{8�.9�ͪ��?9wҩ���M&�]1-n~��9K�bN���sT���3@*'{�|UG�t�i�䴌���|;�TTv�+}o���P/�M��L'������3��La�����)�_)g��d�|��,8�g�g�~��zm[�����V�L�qfC�Ǜ���X�3��I�X]���u�b�R�R8_������`XX� ��oa�#�ؒ�fڈ�0�@�kJ"|&�W¦D�bUl�Fi�#:��cѠ��}�p!�p`���d �9eڬ�b��CLڎ���[�����K0�}([��!f�QRe%�M�|K�Y�Bō�T�"�	m�xf���|V�y!0��/���+��+ ��@Iz9��#�&�����yG��`jyhZ�?+&��g%���������.u.�I4]ł	�<�ܽ�l���}ȡZ?�1�֩����r��(���y+z��L���>��y4o�j�^%Hрކ��:�@o���p���?im��_�E6KW'u�2�N"|'���D��k$7��
e� ��D�@��ĵ��uLQ��0�m��7S�I��IZ���!���4�/<@E~Մ�M1@3=tH��?�6s>H��}�ӭ���j��v�8�{5y(b`�|���_R�XO���GӷxmT�?�X^�!�hMĉ|��]\�0�yY$�B�Z��WA��B��/��{v�����57so��@߆�v)����c�wm0�B���{Vu�a�«�k��zWU��4{Q�1oJX�`Lay���Z�.�N��x��=C�_�̍b��zr��!JޠСFE��ZS�;����aM�]��@�}U^����F�Ť���c� J�o��w="�ܤ���ˌ���۸U����! /���*IL��`���QJpH������ �����c��Y?��K�E=�v	^g�R��҉��=XA�<�<ƞ�1I��i��Cv� �P�]1@�{Y��dJ�y�-)ễM�ܞ���z/��mx(3U|e���Å����z��f�٪T�(321ޠ_BT7��4�Z+� ������mR/�@ ���a �V�k�F=&0��ê6�;�Xt���?j��I�,c7qA�������0DZ+�m�(��`N�1Ԡ-��M���B�r_f�1��3;���
�-:ھBb���i���g��@�����y)bw��Gx=��<��A�?]{�ʱ��Dxt%B{���Ļ�S�D��?��/W����G,ͱíB]�s��[ނu$���QM2���Gb�]_���I���"I�,��Ș� �������1u���}'F�5ˁ��q��#m�u\�d��a~ �lE��!��l�_V?�4>/�QuÓ���E�)�E�4O˘���{����P5;&�W��сA�fDF�b%5gG@��e�\�H,q�-{?-S��Q�����O��L�^�Rl�f�8+�p��!�W_`� ��t>4�*��̤�oH({X�ZqOLv��������J���X+z�vI��D�7 Qz���U���~�>y\_(��=2QXkVf7�_	�qU���bJ�P�i�ց��(��I��c'5������k��L��n���O�g���3U��u���D0�'�kK"߄�y�٭?Mp�؇�>L�h&3+J��+����ʣ�f�P�)�U�V��	�㏥Q�Q�f@m���"HQڨ�f�μ��[�]�D~i������6�]X2X���ݓ��>��
���߭Ml���|2aZ#%f̪[��hQF~��.�I��46e�e�x�NN�]2���Ħ�I�+n�������!��u ��Tsױq��P�Ї��C{�h?��4�Q�[��S1SK�z�����>�
1|pr8&�����!���q//�䂗O�%�2��-O���3V�0U��7W���M�FD�$���a���8˼��z�9���-�1�n{�;پs��@g�/��j��������'l=!+������Uᑏ,"����Ĕ^\�Y�c��8ں�»]���@#ԻN�ٱ��Tc�<�����d�W!	�O�_����8Pq����]w�����TP���Y��T�=+�]���Ŝ}���+ �
p���t&��x\E ��o��6��49|n��i�ۓ"9\6�	��o����-`oķ��u�U��y`]R���+��s��M�3�ݶ�b�Fh��b�i��Z�#WK��p�L�T�c1�ؐݟ�%
�cFW�y�Q�2r"ƾ#9�pȋ�V\D��� b�i�f��nK�b�[ ���;쪸�C�:ne!D˨!،��r�J��<֬�0�(�j{]���g�Q�E�=C6� �s���Ԙ6���<��d'2ъj,S�Oo�ػE���u�b��fip�[�KbD�GۇNxO����ź��RZ(O�Y[���c�t<
Cm����Ȇ��S����	(-�dÕI��{�P���r���C
�v!�J�9V����T�F����L�Z�o>(����`)N���~�[�"�=�Y�d�m|�G0;�=������83#n탟���K�2N@�����`ӝ�-�����.>��D�:�Ȧ ����|v
��@Xc��c��3�`� ��7��o��ύ��:Λx$o�pȠ��v�4�!�W.��5�RE1���]oD4t����3o��xX�����d'���@��6��������śK*��ǻ
�4�#��9�CS|�Խ.T�����DX���s�7��N��͡-*ih�S��zbq��{6�m��[�Oi�\/C�9���j
�{���k�|�S��I53�F�(��ȓq%��!>س°Y�-[�~�v��s��#:?���A���a	(�{�@?�k�ߊN
���I)���þV�i�G��͟$��c�����r�W�����&��?57ޙW��q��"T�������c�+;F�/���l,�A���� ��ܔ/�5TE��?A�J�l��c鐾r� �)��ί����N��a-�����9�4�����!)a�/A�E ��o�h>'ی4���
�*(��<%� ����u3�i�gȺ�{�?���C�Q�1Hc���őƘї-�+g�sRM����_WFU��h��.�L]�mCE�!L���PR�7��o~w<�X��m!=�˥o:3�C�yT'�-�������a����G�BU������%K���-GRU�iKxG+qMݕ��J>�l����Y�-(�>f4���?�3�B�iX��P��X��,0���>�mzhO�S��]��M�sʅ}�����m��P���q��g�[ے'������KL�O2-��\���X�����;�V%d�N��ZfIS�� GZ���xV:�^#&���|@�(U�*莥ڍ�`��>-���C���-
�9p���x��!�n;�=�����������H���C�z��IhxY���,� K�ڇhx��c��/�u��)��W��W�sU)6�G�8��V���$mA��:��ƻ����n���GX#�GcCe��E�d�<�1u�f��d:��l�kj��T�SZ���5�+�?��TQ{��lk(����HWi�w�Ga�S�<�I��O`W�paH3I��',�͚</2�����ѝn���M�TW��gh%���|�\��`c}�a/fE���+����ˇv�#/l{_x������&Y�����ޔ�	5��6��mR��aڇ~������"PB_�Mg�~9�鐍B�d a�~٧��\�������oC�U��E�;]���? �"�>���;�j���/������
�n��x�jM\:�x� �6���Z��U��='�b�*~�:�#S��i
ǁf�[���ڙ�_�?����n;	ç�\Z����x�Ƅ�tE]U=�"���{a���  |��T�Yd�,�.f��[�����*����dB�� b��\NFi�]�Z�#��>��o�k�/�mA�	 b�8Hwn�_=T�f\�
��>�*�ו����Vt0��5�6%	��Dn�WQ*m������O��s��?����d�u�q�Gׅ ��w�_@[
><#@���
<������C	Y�=�<�U0�m>��X�X��qG�b[��]3�%6Ҹ���^�U�*��')k�ro>|��-;�Hd�Ye?"�=E�߮��h�W�廊n}��e��%��y�O�C=!;x��}�u��<�=�i���!)$��)Z>�,{݈Ol!4O�X�`��x�0gc����/�  ���&B���/��O��i&�{s�i!2J�^�?��Nw�^">i؎҉�b؉����b׼����B}����?���V�75�J&�](���D�H9�}@q�_J�j^�������.�w��@�V	���AK�h��`4۵&}�*7��>����oAd%o�,t2R�c|¡�V�y�sAK1�LG/��cѤ�j^&��d*�p� l��� �����jn@t�:Ձ!�7�I�t<����B�=��G�udQ
�񼤏[�h�1���:E�S?�s�P���|�k'z>��z�G��_��^�5Y�"���͐����?܌�U.����37\r.�V�}��������_��LݲF��D�������Q=1y�Ϫ�|���HE��aE�cġ�٘Y�F�?ۈ��)�!��`<$��á��{Gt��i���+�a􌔏}����7`��rAU��Y���V�D�HB� �w;ㅢw�6�2+�S*�m-<��I�vՕ�nhJ���Ͼ�
4
��Xɱ˺n���l�쑌¤��	�=���e9>����$t�R>Ҙ�)�o�G3Qv1��,I��5��^��M�x�P���agu��U2B�GV�J�k���#�l2����������*u�W}�Oy�j�m�����f���C�Mˬ0����"��_7zl���4��>�f����l��l��6"w�)�o�8Vv�Au��d)��F�	�X�Bsl�%��fujM/�0Q?�<h�io���p<Զ���"�"��>L
"��*A��8h$��g�1��O�i){�E"׈a?��h��]4΄hR�&N�C&Pl�1���
Mc�\��'A�=7�[�q�ݏ�$rT��e�~:�9�~��7�,Z��d�Dz����J)[�٣�
�2?F�yp\~9�a�&�w���>�hq�`�_Ϭ=u���z�j²�2|Kt�w7��\紸��#��]{Qr+�jo/�,��;n�óh笈p�a���ԩ7|���²�87.�a��!�:g�wN��J���g�\	+Ӑ�|qvoD���e�q5���EM7�TIJ��{A�#�J���^�?H�a&m�V��w�[�g]��XO��
An	�V)gx1�j;���C� ���]C\J��N��j�MW�T6w��:G�����`�P|�M���i��D�#uGؼ�x�����nF�6� ���8vp�-b�>+�Bu�]�-�����Г3��x�x���2��(������w�����Q9��K,Ǯ��r\������<^ӟ!������̈́=|}���p������#^���2D���+X�<Y}����%��U��6�{�aV�͎�J���Ya&��q�!�'���N:w���@��&�H�*�Z4]*\�J%Q-8b��S��b[��������,�r��fJ%o҈�c�\�=PyJE?�9��uށ	�g��kJi{�fއ8�<��[l�r���</�>2��L�׮`�rl#<��r��?R
Q�#�C�j<�:�r�!��H���4�\��D�D-.C���L	��K��k�ցU������3F~(hw	":�;e��Vft��Oיlq0�_�%��{�V�Q�?"�2���`Z����i�孕�����m��S ���B��ǫ�ӿIҤ�Ul^#5:a�{)uD�w��1.1{%x?
tZR�g���XwM�2�6t�">D�{���Ht��Z���+
8.�z<B�s�Xa�'9�}5�&� I�$OvCsV؈����f)(�ʡ�PV����e����E55�I���ل_�?�,���A�qx*r�xJ$pQ�m��� �%����I-;�@����?"o�I].��B��Q�jb<���1
؞u�5�p���ȡ9�M��Mb��s�V���7��;�fs��e%&'�_����C�ǾF	�eϴ;v"{�Iԙ�����d��R�9e��7IIwI�m7*��g���q��p~u����\���$���~.�6Fѵ}��uj$��9�{"���
���E���d��]J�L�xEW���U3�Mf�K�?��s�@?:�s_��N\��Y���6^�_	�v�6��~ii��t�.�BB��?��� ��o%�~�JG$�9&�Qo��k��1y/얐�p� 9>kۊaiC��06Ȳ�ҡ�p��T��i����$Ђ�$
�/+�K
�~`�}̐����� �,j�P5�x�A�_Į�|�ʩֶ '��4.)z�1nK��. =�����|��<��O��L�L�*I��Y�'�玔��K����o��E�M���R7HW�Tu_���<�!�s���v��L!/l-�R	g9��p�?���h���+2�V����&��T���;�ar�>���J�'.��V�	�4y3�%�S� KG̎�ţ�M������U F��w���hf�Yc*���7��k`6и�F�@�/����ą�1��	�I���٪v����a�����9x��/����~��[�MhO�:<648lY�y�k����Q�!Y}�y'��,����\�/�2�C�g�|�"kFAK�6-n�{%Fl��w������P�kz�e�Fg1���v�ϡ�YS��C�A�8���Rj)�n�ޟz��/X.�[�(�39�jh�L�N��L��B_��>��p{ֵv�G��.˲�*��FD��`�:3���V���/�=��~0��	h����;�r���O��5-�㔛�K�S��U��v�ͥ�e�$��ĭ�0ʟ��Y��DA��-�%8u��^E�I���!̟�+�2k;�������x�m�Ѐdr�_Wٵ�O��Qe��]�)�F&jSF�����1O�AӀ�ጧh�
xXIW��UP���Yۛo>v<�LчBh�vZ���p歂��2U|Õ�yam�(ox5�[c!�tLU�ȫ��sU�d��������ZOیt<lW��d���$i��쯽Y��ɗ�1Ky���9b�T'�Ki6 ��R ��fRI��۝��r��vi��)H�@<�` ��*�썱č}��t��(;�e?��$g�����{�1�������
BO|Ol����鳙	������I%�"��D�4���W�1��71ފ�ᝃ���3\�RP�P3H$����l�[ _y�Wfb�P��`��ؘ�y���l��;��}V�k�Ҭ.W��,.���� "�a���Jh�<4)EK@��N:F�I�:��۽��W���<%_�!�o6���-]��Ц�*au�$�8Q{�D���6���S�Uk�sH]�b�g�~�]�([y䯟m)H1T���T+�m��i��6�Y��0��$c�%�i o^n$!D80F"���Nb����K.�Tk_�P"9��>��6�T�0~���P����-�f��xg��Om�㇥;����(}���-G�Ӫ�S�R0���0��$�]Ҷ��$��Z�������rZ�ZJ��IA� ��������tfsʴ!�S�s�YX���b�=R%�4&��^��BNWN��<W��v��1KGMx/9�G�G�wO���I�e�F���j�׹�WV%��z���:�aiS�l��3í�L�'&
�uը���S��K��D���x�����V�L��î߲3>I���Fx+��N�lhH��S*���Wt�s�i���{�P��L쁀��R�h��{�>Dj��7����!,�Jz��.Ǥ"_�A1N���X���4�����8Þ�y���')�__���#��`!�dX�X��l]Ƌ�g�˾s�~j�����^o��@<��F�Ja��Pz��m��e7�_.��@r��Խ.�~3���¨Պ�j��Fy5���R N�R�0����݊�����+�HՍ+y_2+-��z."�6x�B?bH�M��O�[�O��,8;2,3�Ɣl��������oĸ��������?;.��@
E6+@�q�'OJ��C��`�n){�2&��φO����->�8{��nK�~��'��Ϩ�o��%����I�~h"�p\:8u�F����eQƉ��O��4���Ps��T\4����5Ƒ��XG@K�E��7�9/g7�& ���b]��1�� k��uh���A-fPe!���T���#�?#�9�Ђ���3�^��H}J]�ᄼ���5	�0��y��絜Ֆ��Lg�W�\�X�-xȈ6N��������7������N�4�/T�O�X�TJ�Rn}�ӻXU$(����5z�N�ߌ7n\jnq�U��X,��Ʒv�����-=xN��!����ebB0kS��ֳ�D�Q���F�?H����F��x���e�wH֔)M��bP��ܭۿ�d���q�6o���c��X�9QbsI�Yʄ�ЦV���$��L����݈�j��ŗ9�Ų�E�Z��7�7��(�h>�7�f��f��j"����m�]�/�:vv��\Y��Ͻi�4?W����G�'�խ	�~�	9\m<�M�GC�O�bͲ�����U"	����ׇ�w>�ꊩ���8 �>�ل��uξ��ܕ�����љٛ�F��J�K��U�~���0�g�c=P��f�>w�D����i7;֏"��ΘEd��*u��)�[��D�⺆���y���7��h�:|�L�B����{���85�f6���¹�.�ƪݾ�֔2+؏zB�J��p��evX�D6��v�d�+g�?�� ���(fe+"�A��(g<z��mm$�K(���� =��d��ʙ��O��%G��kM��xs8ª�<���t��VD)��[����e�B�YӴu~=-a�ԏ8g���*���N��a�N󦸊a�^��ˉ�{��3g6
Z�iAۓ��ؐ�����WZ��pM:�	� ��I��XK抆��]�\;��(ԇrl0w�������1z�:�=�	����!�8�,�q�L�o���M���UǂuHT�A�r4��H� A�<ٮ�4>k�
"@����=�Q��Sx�h��D Y����6�}�7�*��$GZۤ��Q�aI��o6��h�)�4-^�u�%��p�	���-�O����y�Y@�9��y�H Qv���&)7
�m��8�ٷ����q)Ѵ�/m8g�3�qC�?�)��щz�sr*9���հr�S�M�&�!<$�"��^���)������N�*k@I
��J��9�`�������5t �®a��o��~o��]@�%��'b�8���-����(�����dp��-t�s��o��F���5'In�Kg��x9�| ��I�.v
�3Z"F��Gx��p��6j{t)���}�_����N��<�U��K�����x� I=�r>��b��E�Q�& H6q.�:��L-����-�����U��������5Nct��f���xB��r��h^�kN@F'�T팲����Zr`?_������V��Ce��(T_��O�W�ꂒ	�����'c�()T��ȋ௥[nx��܇����_9FH�"E���������rpۑV>��,�Ow����a��OqFCaM���0q�"w�_��R��a�r�F�Y�^<�� x�`p��X�/Ζ=�A.4���H�����T�FW���bD))�H�/��*�.%i�%`���5CG˄�}M1z?��q�Dݹ�=@h��z'8�߂�����T�L�Zi���5I:���Qi�L���U���q��4�s r�1��?���ު�p��b2�����!}F�:W���F�rϹ�L���������S� v\q# �߂��o��%���EOu�G�Jܔ*������H�y<4$��/��2���gP��2~MjOR�6%�%]g�'
p_<o�<�7���l��0����>d �:>J��y�柖���e�*�E��\}�D��<m ��{��������^P8��+xQ &Y8����G2����f�Sp�Z��ލ��6���
�N�|��D�LE�6E�p���c}8��l��L�d�)��?�4����	'�xr����Q�@r�U�*���,bw4/3��
9Vaf�s�9ڂk���=*Bu���@x�J�*8:ԛR��ŝ�D����=2���s����1���KWch�����@��e������sq}D'����#*�g�.�~���)He�i�|����|ӗ�>Ҏ����F�m|�u.-�y=�$�����k�76��#l=�iK�n��ꯄ7�7��m�7}�#�;��~�2ZR_�;�<�`� ����&�T�.|&�������o�T:�'�ݷ�ۀ��[�%�[��?gG?P�o i�J_+��EJ���X���%P2O��(iVh����Fk�'Ob��.s�&��t~��;�˪�E,�@=:={��-?��t|�b����Y�l*B&{]k�\��qu�Jك��``Gy*D(	�Go�� l���z 5[�me�s&y6�[�����U�̒B)�7GňaۦVB�O�S�	�����!(��]g�4�6�k�(凨���ʄ��ݽ��a�q^e"y��S������KwE��]+h���k2�ЪI-�ٕ��x5�e+b\���4��m�I�����-u�g@�@e�	�!Y&����Q�Ƕz�0Z"}Y.f�X8wo�R w�!s��rj����Qe��7���-Z�F}���L��O��U�x�/�� �BM�e�V=�"	o
�@�H�V�'�In3���]o"<D�KSTm?�μ0T�>E`��_^�o����}�ГǺ=M�*E&-Ɨ�P]��GC{������z��q�r��|>[�Cs�0DG�S�ڀ��4�O����&��>;�솸Q��_Vnή�5z��꠮t�����X����z�qAE;�q��)�7��x��	��(y��=7`�Mi�Yo�O��@�X� 8	pL�v��J��>8Ü
�χ!�_�����63��t��_��
Ǌ��O�'��@��F��4���fG��H�ھ�1�l���ZZ�إ�ÿ㌁�,b��a8N]�^q��I.����(U�;���,��Ɠ��ʖ(����!�A&��������h�H� z�dV�Mǜ`Hm�Έ�	��&Ʃ�-�tsj��JϷ<�XUӒ C7��"	W���f��S&M~r���D��^ne��Ưv Y^�]�%�q�?A@Ҷ����U�_�U~��\��r ��(�	9~P�����	n8c
0Y
��g0�ρ<$a�<���ЬeE�� "1�?�k� ʚV����6���>�+��DDO�)7 �|�P�PJ�l{u��I���ac�����1G���1O�񣒾Kk`}0Xm��}P3�da�����.����C�_s�:��w
���J@L��տ#���8�$�,c1�)C�]��A&����b<���vo�	�l�a��G�Y
����%����WB��7��o|Fs��{��a�d�����T-��F��1n��7���?��p\N���(��i�zHcQ�[����=#�v�䮷������j�{���&�}(����,?�E�Y�wY�V���r\��HX��M���c���	�E�T� �!� ����ȉ&��I3C�[&ow`1k9�]��ؖ/[���*��3ig�bg��X�n0"6���(���J�U�6�Λf/�a��
��o���'�����_�JfAg:ۇ���BW�y~_pΙ�0�%�O��oM�� 6�rf{�~���
������{j۸�Je��,یFU�"��\j�3Q%!�;[��?��&4p4��2�_��l�p(���7:|����I��֏���݀*F$�˰-��-�� ��Ӛ2ܠ���ptZlΟ�
���5V��QmM��d��>���D�h<������\�HS���~E؁���J��2#�?�PQ��TH�~�$N�d*�� �5H���.�l�P���,Zx�}Hb\��Tk;�����A��*~�ֆ��q�X�U����Y�J�ej����t�
�jz^�Y$ ��da�7�����{�5���Ѿ�@���э���3U�W��6�!Т��y�)��Y��� �N�3��wo�������2�FC���,a\u��.N�G�A1�ܑ~(RV�|p�?pW�R��p�.nM�l�Ʃ)/�
�Q ���Eo7�L������:ף�"�uCH��x����+��oj���݇�w��?�����c�;Ӱ�G���&٨�K�4f�d?�r���i�}�Y�v���-�u�(��(����zH�:���Ӄ�5L��Ud)c2$G��aK^�tN"�2�-��9w�K'�)�ܢ�m���e����Q P����(����<�Y�{Ȼ.Æ�4҅{��$�����Zp�TWE:|W��WD�7r�
n��6��fv��/��Z$����G�1�j��s��Q*�� EX�0/�����P�e�#�)��v��u��M\ޅKh@�p�2ןo#ٯ�?����p��!s|8/�{�-I-b���rV��Đ+ �ɿE$�4��;Z4.�2�.�X�é[�T������#:�1�o�H��� |Q
�9Iq/}f��Ѧ�(�x˚nSqnA�}��$���{e+_���f=�C���۰`� ��怦�2�^s`a_oq^��όWjp����\v������0� �x�7P"Ͼ��]tߤ�r�E�3u?�R�򲩖��[ج��ۥ�+����5�0�p�g����y�NH����{�d��W������sb��>i�~�:j��¨�*���}��f��7������5� >!K+:'��}�R�J�!w:�[�;F���Z�
�f���[3� ���G����.'���j��0$��}��؅�r�����_r@*��A�m���L��h�:�Q;i���
��6Op�Z�P�a=M.[!pl�ڌ�|��kd0�f�V��	F��
F���iO����L�Y[,:N�m�X�|���L�c���)�v��A���k!e��G=$���o�c�#��3{Fߐ�����ƛDS�7�N�*����T��������Bė80��y[G��1,տڊ��
N�ꫝ��?��j��⋾����E�
)��B,1�J���
`Mʪ8�\(�bQ�t��P��,/��
��-�}μ�_1U����ދ���uêN��|�죤?y�(3�u��s�8x���<h�p��G l��/�G�{��Me�o1�8��Zy.�8rW� ��e�!4",)��J�ŉ��ٕ�4�n��q�7�Gd
��3�_�!�,59�NtN:zقFHJ?C��P�z��P�0}EmT�w?��^� ��V�v�Ì�laE��NK|�wQ���q�8l<��]��.�#TqZ��@A-����O����Q�-O��,�?ҡ�mc�=K���M�a2^bM�o�`Dߤ�����7���w�WI������u5����H7�;ɂ{�@��ɍ�h��<�1a��֠�z<i���#�+p3�˫���J�B�JB�씯�XJ����C�И�=�7ĵ��4��x\�*�X��"����\N|�ؖj��"��tR����"JR6�3+��_r��%�ա�m��}�@�8��"���h����+nJ�PHti�E>�m�rC`�p�q�dj۞��r=�Fr�J�k�	�}?��,I�ضy}�
  �=���W�>_(�ύ�K�����9�i��������zE��`u�*��ms۶�V����n]<͖x�xtɌw�?�[O���ߖ�:@	����}aڀ �� �M�S2Y@���})��d��:�$�w���ȉ�D�
JC�r!�\K���� �c������N3D��lG�6O ��L�-���ٍfK���u\ S�%e�ہFH���?t�`r%��v�{������&��[f�eD�e�k��pdPo��EP���׋B�g �Z�Fj��c����ZgHWC1"y�P��̻�s�SV�K�J�7$7o��V��BdR�͟ݟ"�w�S��,���$���ݩ8���w�������w���S�����z�)���	�a��`_A�U%k�7���Hy_����x�F��������K�i�,yYľ
��4m�nζ�z'�V�x�;��7.��u�M
9� ��c���0P�G��z3��	u�.����j�E�G=�OO>�<�����-����Q�q�;�n��dAʦC���@S����<���� E��X��W�F�
���G3E��<(�[�-�H��p
�DX��3��BLk��6кT�9�o�P�@ű��VkE/+�Q��e�(�^�<
N�h�_Iݖ�,h���	7=��u'��A�'b�Y��;�m:��0"��|���w0�[�f)D�7��,��Su�r���4x���;=��<EiI?��Vw�8�*���Gazh�H9?K��3�/��j�Ęr"ڸ֥I��[���\���i_B���JA�LWp)��-W�<�y*	Q׳���j��]�t��*R�yBv�h9�w�����V*�e�1�tz��٤���d<���OE�����k�3��P���b��?{9Vܥ%�'blˊ�_x��k�W΂����������h:���^��E�k�G�-��hi�gH,��8�P���/�8�r��������C�p��a�{[�Xt����O�D����(T/�h�R����3뵎�~ �Ynt��K�%���	�_��1�n��O9"�*E��u���ۀ>��y �|��q����F��2`�����l�b5�,y�}�gQ��_�Y�@�I�+@���X�fK*���Lc6�V���"sm���Sw����ή� �8_{�VetX��Q�����Cr�1�q�q�b,��#tә�o�8���DJj0���4^���s�'r��z�O�F[2��i}U�h�ιۈ���Q)8�f���ߴ�:g�ڴ�Fh�9�X��q�Z��N��q�Q4�hJ�|p�o��$M��p'���r�-*�Bʚ�O @QX6��OƸ!a�P������de��.K)ZI�_���~�!'�o����2jۙ���jɯro������M���1�����~��ٷ�s���{���ܖ g�9�����t��;��b���Sq'lů�i�O0�5��]�{Y���G�?+�e�����Y6 �cH$����(�r�������+�&���;�*(���7�|�
�|��'�6��g�A���]I=��#)Գ٢h8نȲ�13H	���s�7��s�*�!4w7?{�����:a���@��c$K�,��T���Ct���DX�l�myt��~�%'f ��J���'����{˪R@�ú��{�*�G����Õ�g��Q�p�}�GӖ1���LS�"�rD{=)�@�Rj��^<��/+���G�4�LF4�[QQ<��+8DP�H��z<"F�)m"�7��5�U:���"p6��=���^ċo�v�Q��P��b+��W��l�����-����*�8��"l>G��E�񞋴vPH�r�L��-Z�d�%��a|��������$��n����,w�IY+�$J���w�(nMro�2�Ik��|"����7>8%ګZoϏ�GV�w�.�����1���ٙ����ٗчYȀ��E?�a�֞iC��W��I&,��4ʕ�ג�aFWD1ro!�熃\W�ڸ�/�B��s�T{oiD�㛨	��Y��<� �m�Ľ֦6
���3�Yx�]�$������sX�.oWy8m21+Hl�nUи���'U,8nW�ſVz%oÂ��i��{'K�xg�zey+���+5�^�����n"{��
K�oX�S��O�Ȩ���1[1g�*����^��~Q�%&auO�>��Y�4QnSl{�y�P����$��c���Q�^a,J
}ăP"Vw�{k}1G鄵�Ҳ�����Ӕ�eR��#��U33�yq��z��:4�_��1���	��0�U��ʚ�?Z�X�XP� �Ɋ̜���թ#C��<[�y�IPG�����9X�(	�gͤ��ċ���t��������#�*/��+�m���\��+��n�5r�X��ၞ��0	�!��s	H����"u����[`@'аu�軖��2��g�?�)ұ)E/����16!$�][����lŰ�].�6�}�����I��t��V庂^n+t�`�u`";�,���o�:�e*gu��`lZ����.v��zUKI�N��
��H�"߾��a$RtS������P����\�^k�LAk��G\����"����Jp6!Ϋ���#�%��L��oWpܸ� ��o�F��P[�/
J�S��2�aL;�$���X��8
��?���-2�f�{*67�zŮ�m�@FU��4U�c~˲����p�"����/j�*�$�k>9�"ia�<��T�W�-g�rC���c�d<#��y��>�H��a��sl�T��<{}Ǫd��1�&�ˍ���X�Z�#�:�ƹN��]G�~zx{����K�����������C� �7��9���;'�0+�n6�3sL�An&{�l�nL��,��sA7f��ʍ����� �O���<N�/>;����<7P�ITD]��D���X9fnfP���֩��:�"�]�͏�Π�R+�������)���
��G�]}� s�84[����`����Ѷs�鴲^c��_�������O������J���$5�����|���Ȥ����������N�a�Q�aVQuz��@���Lb���u%E�V��}�w䫖Ȉ���lLln1�D�}ˢu�����D�)1��`F�}���`�Kk��!��'{.�3����H�@'zޞ����kHN�8�����#d���>-%Z������^�j�s��beH�i��Z,�M�/�;_()��J*�����-�@k�C2�y���<���Ԩ_j0ֲCۨ����	���ˈBVZ^H�B �K�3&+����m[b�T�ξ/�Sʚ�z�TZ�̭����x-�ki�,n1�7���[;�W��E]
�ݪݓN3N�Z��&���Yב ��{��Q�}j����+�j�9��s@�W�=��y��d+e��|]�<H����7|�!�xBWQ�Y:��D'��:Ǡ�[����������T��̉RF�-�v�S1��`Q�GYɉ}���~|����:#	e�j7C��:�������YAi�5�j��Tf:��9���;Q�X�̅k���h(X*gA!�5����N��[�|�$�0u�_f��@c��ulY��,_�����9Z��(�~}���c՟l/&qe^Γ�FQϼ�ӟ]m�P�\$DC�Xi��*qc=�ێ���{O����J�9{�ze����Q��,/^���rJ]]�tQi��)D�67�\)J(��s�e)��yI��jZX�SDf��dgD��˧h��qh�gt�:&�����sY� }���!�L�z*HU��;��:�����8�6�|a $�Rc�:�$,���Y��/
��%��R5�O~�����@�(>�����z(��8z4�R��,گtyo�jd��T�դ��2+R��	EM�H�����*�K&�b�n%ԣ���MK�O% *$;4��w�j�����ES-���ؤ��`�IbU��<�b:��;��"{I����쮛θ����U@^�U%GL�_oR˿y�ew�=�H�FF�݆K:8^2��xc/�,g'���I��v�e�����\�^ח�9�t��v���=4�!]�%�ɲ+>���sk��e�+ mL�i%�db�Eøy����kXZ��Ք�63������2ń��N
>�)��PX���F$	��Pf�R�Lb��X�N��O�:GbV��58Fz46���ʓB{�5�L8eW�g�~T��nfT�򟉾��o�e��dz�^� �A�SV�%�(�����d��5��X���HZ�7�� I��J��]�������N1.  ��*��=�n\#���b��~�I�niH�ڥ
g��+�,�
v��D(C�L��]��熔Q.&K|�Vv�^'��X=ؚ\V��@=_^�X����#.5?g��L�(���7YZ@��8ԇ!�i:�EŁc�0�K n%#ݢY.���1��P~m�
���(���l�%���N�H^OurU6�����ڼ��K�=���,b'>�9	�Ua�nsh�h�OC��g���}�}����Ũ�M4��~�fa���m2�4���1�O���M�-I��m�Ȋn׋�ޥ6����ə��[��|۪͆l���K��㱜sL���Ҷ��CL�8;��v�W3�$��F���㾪��i|v'Ar���e���C/��w7|bM h��q�W�ʄ6��/�p����UKX�Yf��m�z�yGvl����(H4\���h_rщ��KpփV��}��[ŚKS,�F�[�r��h�!���d�6���&���-�blU]�y!�	�/:
����}�;���� �Y�(��:�� ��>9�LC�wC��0��"�!١�FΉ~���\N�}g}5��5��g��xh��M�=l�L���,X4�rྛ�-l[��ix%d��w�u4j�5�hjZ��Ւ�w0�����1M��&?�䴥����y̵;)a<���`��>Sě�x%$6���,w���tjAB�~:��n��P�%�	�!$��=1ٶT��5��B��@x�Wݓ����M*۵�_=�`\x���۲�b�ڥ��s]՛���^l�&zh/Q�~�;ߊ}�O����`��;4�Ϝ05���0 w�uK�0
����<�tm�����֘�юō����\�����=�(<P�[T�m��z���{g�5��#��Y*�l ˅g9�>�Ol���²��?��J�>}ɡ<*f=z�ɇU�ܷ���η�v����K��Թ�Y�/'�S1�H��mo~�C��uߟ�쫄�ʍ�(�]�%b���Co'�4Z����*����!�w�������Q����z�_Dv��t����Ц~5Mr*��]/�{��''ɬ�1GΎ�6��	=�K���&X���A;�DyX����WVmw������뜤��E��|���	r{Z<�`��x��������("	�:���5a����L�^�-e���W�g�5����k^��MC��|O(�դ��jje�A}׌�Y�t��Q����A��'�d�]�Q�P�;��>�Pc�G�[����;~�Բ�#b}㴆����� @/�}>��J�ﾭJl�cIls!��зֱsMXQ��`�q�>yW�x?7���S��n�(�����������QAp��<3���� aV�Z�[�	�h�`�s���S>����Ŏ�I%S�#q��ՙL��wh��]V�j�������SAR�Ӄ��h�Ҷ���Ъ3�N�o��*�e�VAq~�;MB�&�Ѕ����p�xu�rjޛ�ѩ�u��x�r�;�s��7����i󅒒�X����8�Ta��~�Wt(k*���sL�$2�'C&�B��p��)4�^Ή@�5�Ф�j��s�۔�ThJ&�d=;bu]Q3�{>�����̝��d#���X�=>�-D2�K�AK
��>y,�)H#6W���]��OF� ^�Z������N���|
Z���V S����s�8?�)u��'�H'� �e��Y�x_k]fdW�8���C}!Ŭ%h�Z��j��]��O3�K� ����*��f�Gd/x�߉�/����M:oD
!ӧ9N?d"i����lg�л����l��M���;�䐁zR�@���m6CI���R�ΐ��DL���y"oS0&�?|n����ۏ�AB5*ҿ��d�.svp�:$����xR��E^�^��S��I{k�����W�f�a3�[G2�(])��*��1�5uR�� ��2�MJ23_OHnʱ V۪��������e��19YC%��������j&P�nID�eit�cń�j�9M�O5�\T��M֖+t	8�L������t}ytG\C�D��E
���Σxd�9����.��� u�X28�F� ���
3�P
VU*�����ٷ���[����P?J�`S��&�d������J�ֶ`K.t��Kʙ�&����ҿ�;����d\)���$�w�I[�9L	��B�Rz��N[��k1H�ָy��RP>8gؿ��]�w~�n_7H��Rh�|�N$rlZ*�a�Hj�NA�`ką�.N$�yy�P�z!����ؾz*w_��E8�9����B���Ny��p�}��hR�� 8e	<�y����q�� ��'��
��5��A���\��zv�PS�I< Z^S�*���S��=p��P�D��f�O+�"��"ӁV��"��6|
��)
$��r���.n>���H���$����1Q�(��P���Q_Ria����|F����q:�<s�C�7�$�\��6��DJ���)�gH�$ݲ`Yӻ��_�/�QW����ty��+@T��	��(g�u`��ěl�����n��:0
�C"xD3�s1ɮ���KK�^g��fB6�(��vp~���<n?����x�~0�������,�b�v6�8���D��>S���{
��<I�9� Tg��
*��*�U�SN���(�R�Vho�=Z����R�v6AG�+�Tޞ��Rbך�*�<w�P������[ al%��t�	)d0�i�g1M-CS�Dg�� ������@m;;�b+�5�1����b�7�V-�YA\�d��-���f�.��cy��B��oF� g�"q^:/W�yz�k�\im��3$��$������d|Ɨ<+l��a�+��}!�?t`��xEb���u�p%�!wDHv�2Km�u�R�vj7a][M?��[-Ц ��8�CC���ds��������&������F����jZ}��F��ݫD�ԍ����j�r���*�IѨw0[��t�QI��Rf�r�Af�,�6��=�r� ��a��i�N�3s>�E+_�bzn0����r�Wb��޽��x�;�����"f�A�@e{��n�/�?n��i�����	�豎����n��'nC��e�E�6��[��+F���LL���� �1T�xYP��q�q�V�쓃k��5w3���+j J����px��nF��b�w9^l6Ș열P>�x��)����d��e@H^}��4�I��ہR-����վ��OH�{OArtx�����e����S������@G6絊��%��x�hG����;�1$|����G(gˁI�M�6p8y�K,e\�?���,�"6ٞ�Qx�c�ɒ@5f֤0�tV%>�Z-ངmw�l`����!v_����o��`�;Ja~�t���]��ߚ�7���4�x|7�O�8����H@Q�6�CI�D�zKT�{ae!�K�֢hO�w�(�:����";Vvz��@ni,��XSB��ޱ��J6{T?'�ȝ'�DbwN�3����?�<+���e�L[qAlN�X2/�I�_��4ڏI:ZM��[ۆ�(���E-'���U:�R�.���w�����������9kqܝ0E��}��Uy�a��{�S���ǠI��:υ���Ī)��g]I�4�HY,�m�ߝ6#���O��չ�U�e����U�a�kГv����� ��z���)����^�pu���	)\J�I�z�Pr�G�W,űRL"��������4�����f���;���j:��Fl
b$��X���:���F�9Ї-S�n9�ޏ�6;���D�t �`(��\�mD��p���fl���_}���y 8\&x��Ua%�UG�2�̥��Ւ�`��p��%$�&B�I�J�9.>ϗ8��3J��&���f�7@�C�8����`}L���z�چ�b܅�6�J�ia&�'(�P�1�"f�w��M���R�����t�@�K/nxK�H+I?ݣ���&����{l@/^n�=p���BQe��:��O4"Z���C�3-�+��l���-��,$���yj����F���cwD��5�7@��+��Y�J�A�50���9]c�P���[��J'-7�z���TüO��zY�^)u�ƅtN58eN�Y�XxPQ���Ț��>��﫰a�2����$�Q��⳧~�#Y���aŢm�F�zJ�ދO1L!1lq�ӎ�;Y-��������?Qኟ�l��[��S�sn�j�݋e�Tu�����=���n�GN�uT"(�ݝ�:R����M�9 m�L�ڽ���k#�I���@*��Ȋ���-��5�+����i���0&��:��9a<���%��=J-M�������iI��3h`�:��x��Y�`�NɌG�k<>�VV8�@s�(c�q��D0t����_�hZ��g#~�?�vF	��hp���@�]�mP\P�	��B�*g�hk^���QW���7�Sj*P�X�Pl/C�S�L'�_�m:�Ǻ)��?����g�r|�!�9�e�0'��Zn�B���=9Id�r�&,�~c&��F�s�$!P�I��4m���ܯ�B�AI�?پj5�ϣ��������6�I3�!K������U��#�s�;:PV����Y�3苴���+��-؏T3���U���,��y��v�I�[u�h��Q�F�w�+��?k����&�i��C���9Ad3��N�ǰ�4��6DC�V�Hk����J>��af(� �g�5~���{�#�xq%�%൦.��a9� 1��͡�V��wX��o��1C7"#*��:�<�V�����n�䏥�ê�zFg�S �l�U|�:�a�ﻐ���V��9���`u8��O�T\�]�E��'1�����bY�F�	L����5�Txvj��F�΅����A�!G�<����yd�_�<��:�����^4X&������g����5\����N	yX�[(&�a�3?@r:�Pgx;���)��i�O��𒽲�����n˱�4��Aw��+�����a?tڟ5�>����ͽ�P[z�CXO���p��/.�r>�z35�Β6!��{H��+9�:'%���0(���P�@�:k�Q&�Lj�@��kx�9�^]
˨�* �L5-� ���U<Բ{�s	F��!�wIP�|�dG�_�+�}}"0�����e3�3�<'����=ȇ��j��m�T5\|nX&���]�o����jn]1ta�:��d)�2�k-N��⡇�������ߛw�tQ8��>d��ՙP�/�S�K���Q��;��z�8���;2A���<JK�Gg�rԝ��qeNT�DjTu��|!T����	���� ���%�dPj>M�/˭����[
+�b�;Y,z�wū�ͯ�������J+���Γm��ִ�m�B�����:*�U�-������d˺=�v�I���c��:$�삑���-�3�W;�K��=y���d+�ٌ�uX���J�&'��v�!k�yƎ��Q����;�DG�Wn8̨���Ҿ��u�N4��H6��}����-�;
_�Ƚ�U�R�mmj����6Ѥ�D ���`�О�:�^�{�#[��s+-��N�Q�7�*���9�Mz�)���UR!r��l�Y��S��+���]z�����\[��찟6���%���׿�Xh�F��:���XAW�ߚWk��6ɞ���^���@�]�py��͈���^_�e�Gn�Z� x�x�nm��B�uU`:D0��eƪky9��N�~r���ۜ�~"�\���Y���o���qJs�6\��?F�!�x_޾ql;a���j>��&� �	���Z:�b�^H�]п���Y7 ��n��Yꪞ��bֳ������4�q]�f�O�[wt�{f�`hU�r4^
�TX�9��	�h)�/@Z��2�}���%���Y��lz'x���f`�s>��/�4[�e��0�ܿ,�S`�� C��Z� /��Y�.
��e5���&��ֻ��C�i����T�O�=�>s��oS���*.N(�XH�k�7"�E�K2�/��\5A-r��sw��@����3�FڼR����ھ�o���q`���O6�����_�P7��1	رMGEvJh�v�4����}�������?C^�qוxahA��PL���.{V�����ES@�P���[�e��<��h�w�ǯ�)�a+%Op�5�ϥ}�wT�Y�F�����7���ޕ���k;��K�N[�l��|Z[_t�z/��cm��
�_u4�t�uN���PIJ���sǅ&62�w�I�����@�i�"�B�-���F�E
FZvHaXC	���:Ҩƫ�z
�!@�l���4]Q�K4����h/�h�ρ�i����{�u��N(1$���d�_��r�Į&�>���C��	\�-� KY��|ʗX��veP��Y���!���W����+$��5`�������2jl�tbɏ��t�Cee��2���l(.2	{g�3�Q(�ޓ��W��̑���c�uE1�Q�|>bHs��� �No�$�dC#��oe�o����-��~\��دVy��.���5�7��q/�N 0����t�H�/�"j�]1��|@�.sl�h���0)�'����,�8�s� .��kAYX|�t(`o���%�ح�y5g~w m�a�SΓ9�%���-��o�D{Al��5c��t��9�Ϥs��r�<��D�V�?��Ʃ��r /�4��V"���P�(��!��9Q{��fp� *�
��� �H0����Y�z�hv�q4��;T�.��W����Zhd�t��68��7d�~F�U@|���8�?~�2�B�d��{B����]Yr�p���:4A'���=�O��[��Q��d�5!�,vJL���}rJ�#1�>�����+X���܆:a����ۜ�L����r?+���ev�ա$ްb�ׁ����Ը�($�=�����F��Η@t66��Y��,�I�dj���N�dqSKI���cgEy���x�ufy$k�7"���룟`��p��!� �E�ZW!�1$�]dA逘��aDi AG�ׇs&����`w ���8�5���W�(�ĺ.�K{����]5:�ϖ&	J H���$��k:д��Ԅ�kz�s���w�,��M�&�U��}6�mZ�v�̮�{����-�3�j��"XWW��5ZM�<�_6t\�W��Du�@g2ψ�v�N���6�CN�x��L%�=H;Qa��| 8�Kʈ�v�6x!Zՙ�Lc=,�u]p1)s�^��ʣ��zs%i4
g���Þ��h�=�@��&��F�y�o!v�|������C8��'�-y����0���tt�s{Ls	�!��?�_�1J�7Z{�jl�-`t��M��M�8'4��ڙ��:5�?<�'ZCʵq{��~	��~�'tɛ8���V���>K�줅�ј��Yqxt���㴑N���<�%@����$�	��|���gn����3:�������YQ�]������w�`dF�٣`�uå��PT0x��3-x*�����"�����7z���!5BH=��Nx��V��k���ړt7.Q��%��%��%!��	���>��"x �P�N���vț#�w,$S֖�[n\L�*e?s zc&=FF�ڮ+d���"����Y����[��o|Φ������3�[�~�uc6���6ܹ%�$9��2�"��cHc�xA�{�@�,Q�4W��RB�c���$��E��j��D1^��F5h����y��zX�5<;�cς��5�b�`SY��<�.9��UW����1>!�g�L��9#��o�F�Y��+��pM��$��.&��r���O[a�㱥���5Z<��V�R�iă�^�(�D����}�R��{h��*@�e4&�^q)��?���L��%�D�ml^�5��Y�����+� �'D��\�}!*3� �.ә��,�e��'�M��Gq��Rw�'���^`�Y6��FS��<�v�Ġ�í��N��*��٭��}r:��\�b<}YJqY��,t�lIݿ
��!ğ�2�@&,����~���v�3�� 5���Ꝋ^U�=�E;d��v���Gl��;���1��b�u*Խ�cW���+9m�-6�\k2�VK�l�/����\��fi�Щ�ԧ���x��ŕ���q0��#���f,Ig!v�@�8iH����\�����r5p��jҽ��޵�ga��ѫ�1;W��P�`��Z��i�*%���t�ʘ�ŻiӾ�B�c�_����I�:��rVOOp*>	�Q��T����ka�Q 2�X򶵗�,ؗ�zH�s��]d�-.�h��<�X*j�7�0!ʇ�I��r*� ��%m�7/10�j�P@�`��|��ÒP�h�ڊ��O���'J��GKU�1��F�x�j�xWD��C����g�ly�ɉ"P fP�q0P���x��& ����@@WȠ੆~bZ1�^	�Ȑ��3�g4+�)�v��0iz�D�A����,x>�4��z��+3��з��0�����K ��߾���zp:8l�D #%<�ӂ������d�L����x�2&�|����UM�D�բL^s���NҔ�C1p}#��3��JN
T�ʹ�"_"K�6�w�P9f?����{��q^��+F�EJG�>#��-�'I��Q��i�з-"ҼEZHٛ�2b����z�f�J�+`���fR:95U?\[���^4yEj�Qu3٩�������	A�A���d�+����y�l(��M�hp㱺�������ɊߩD��J���G$� J�~<t+J,��U=U�N����j��6|�'�o�B�����hJ;;k�� ��h���q����ҁ�[G��3�^f�x&�I��Dm��d�]���/���1����tR��4��|���{>�J�U�Itk�bМS|�:��Vr7`'�?zeeW�zw�$Ͱ���[^1E�A������o�`�S�^�ԫ��d)����29���/��4X��~&���Ѹ�ښ��9�;����9��A�5���m�,-"�r��J��u�F]d��RǸ��oE��dG��!A�I`�C����Je�.[?�ø:ԅ"ϫ-!�3��ՠ��nE�78�{H�͹�+��5��C&�Enb#%P*0Rq��2�X�T�Ђ�!vw���CU��ay�_בc.w�����x$E�ݘ�ag��%|��V���� U0`N�0���x�����tAȸL�q��k�B��s( �P����:�DM�iȬ����`�;��4�0��'�_�!x*�2sz������T:=n��$���-�`݋����������_o�4�

{��m_�&v�ml8��
�X't�� ��I�D��X<��t�����(+c���ɾ�����$�siD�PY{3[��XU��r�ќ����P�AFߜH�J5$`Ŷ<���F��u/_S�,�a!�'!�#�{��=%�g�}�3����x��e`_�pb-B�p�w�3F�橢�����|y1q��}4u�Q�/�ް�k
�u���7_�]dO�8���R��UF�p{�Ty��{fg:��������y�}��4��V۲��V?�s���>��j��J��h�rV�d�Z$�Ujgc*��Mdw�$k7�@8��G�`_ޅ?R~���!\��2z�L���W$��˕.nY�_��coS�x�C욞)�t��輟�:���/0*�]KO+�R/�h	ǘ~�.W񃤐�Ĝ��j���9
�6 ����>Hń�	��`+ngMAQ	�!i�0��`قo������E)�(��g]J�q�^Q���TOk���P0Ε�|����V԰8U.YN�y��^���T�Hl)�q�=�O�-�5�]
$���6��"��'�"%��%�g��֣��'�x�ML���]�O\��Tbk�!ˀ|�"�O����g��N.�H�����g3�r�)"�ʺ[PI���q��7�S���q���.O��$��Iْ��S$�.����uvl��K�4�ʥQ9	]\�ǫ�7�׶f�ɋ��BV_m>]>���ĩ��
�|���i��^=�A���<��0l����xu���Y2�*б�����������5��6�6�Lz����l�-T�j��V��R�D=��u��T��<槦�����.%=aI��p��n�Sp�$}�Է���H��.��W�{���Y7�g�X�'�a~�M�����������@�eG/���a���I�1�����p�wؤ�4���I�u]Fᣗ��P���v�8��7���'���:�d q�y
�8��� nM:���"��Țy�6��a���-�F}Я�+ś�h�`Zd��c�hO�!ѭ,/���j�ߓ��B�lz�q�Φz���L�{���E��_�^���BI���ϴ�n ������$
r�u��s��*^̘y�J����4�����.1�=�l��Ԩ7.�C I�%f�r���Q:�Ʃ.��tk�Pq��Q{g[<z,|��5���6��O�G����k��cq��"�����ʇD!eJ����W5��u�+�^ 蟫��>�7Q.��L���&On���l���V�v�:B���� g�HRx��z�[���+��Ns���nH��Z�ܤ$�9+�vD�1ܳ��Mҵ�7:-��������hq��%2 �:��'R�$�;$�d���&�*jnK�=�� c�����.7i��r`E�M���i�`F^P�Uw�{$���V���/�K�e}�82�����ÿ��S��6����	[;'���Q��|���[����Q`Hc�H�nj�Ç�h\�h�+�D�ۂ(�Y7w�0��m�v��=��
��ҕ7�Z�ʂ����lqo��w��l�s��%^(|�HD����J���4yJ���?�U�j���?U\��';���6���/DBpko���z��f�$;���3ZU�i�D�Ğ����L�A�v��,�� �^T.�'�E�����[����� \�ӭ:9b%^��$4�3�j�
T2�[��{�����T>Ť�~��5)���g���0�N�jX�'�u�W)�ob\��_`�vq�<8@ī��}EM��MG܈w#��5r�ǃ�LS��u3�?�z	1cB�zφ)?�^����e���k]3���7JwI:(��ʥ��Z��iF2��}�ռ��=|U���V��6��5�$������?�'7@��I�w�M��[��M�^dÊƎ�q��h罾�7 �^���Z�E!���{�\�Bg+5 L��ɜjد�CЇB��W^~�����o����T���L&�
X��
dZӳ�����pM�f(��WȘ�Ư���^Mz��n(W����4�ʚA�[%b����r�>] 4Iߜ��Z�OU*����hxN>�z�^��v-�έX- iڔ/.��|�g���֗[��aY����@�}Y�Wq08	���#i���,�s���[����j�`����<�y�����|4r�|���%��:���3�ej�����L�.�x������O��1�̠:����;_>��\9O����P'��#^��L�N�&�-��oן[ԡ���'.^��>L��B��L�@@�"����l��f��%רu��W�I���Asac��h�Y}�`�d���-#�`�:��o��.�����:�����d��c^��-���Khפ��P�D��l�� s�F3bX�87��l=m�fͶ����-U����&�%�n��4�&�Ol�ކwXl��fs�*.m��q��/��� 8���)�t	S���S��\��;hJз7����i]T�c�zlž��h���)Mi��+����K���	�>C��w �l����n��ղDF恳To�O{,�PѠ���B�+J{oX`@�HY T�6uQ��)���P�=7�"V�z&g�捜ϩ�Ƿ��4�P�,�g���P('�-0q����B�i�R�83�F���{{��x'�Pu��5�hO����H��K���{�{D�(g�$t�p�}�gM�G or�k����&25��O�	cӄ=C"qk
mo ��,��*o�r�����÷o�k{ϫ������(p�%��=��ZC"V�R��p��	^���8�a�~A�ѹ�R��((s[*%M�#duL>E9O�$�{x5P	XԑNQ��T����]]z��sD*�>A�����/Q��̪����0Sy0�$�2>���$��|7��]��z&����Q����(-a��͸�U���F3�F=��*
	e[4�'���$J8�uI�c�RRS�����p�'{�0���H�QZZ_\N:^���٨�ڷ�n�т��5у��p��30����4�J��=AA�6)b
�5�n$ʞx�3%։weYQ���J��ǓGT�P%���0�����+�4�Xy�`��-���h���ƕ ���\��\у%��>I�ށxk�2/x�t5��I���A' "	9/a� 1/�W4�޲�q@4���_ȓ��1��;���T\T�h����}w�r+,}�6`<�&,�2q^�5�$~�<dSƠ�����}�����/`��W�-1��o�t��� ���}��F��g<�,M���zq��QMQJl"�7@��+�M��>?���v�7����zT(R-ȣ�sy'�|:��<�V$-�j3�2{F��s��{���๋+�@���%���8������w���mr ��t�������$���ݶ��]|=�_���F�!.x�W0��;&���ִC&8A�"?r#�q����a�?�J�b�
�)k��58s޿wER�]U��\S���~k���x���w6���T%2z�3������Vh���]24�e�3�4=j��z#Pbs�c��lj��"\Ifb:�B�[��
�ipW@��FA�E�b�F_6kj=8���4h��])�,�]SD������S>� jv�^�#��[C�}�AùY�����N���KE���eI�Y�����P�lW��B!UD��}I��$� �Cz�Ćo43H��Fl�}���a��WH�!�7�9y"�J/�x�)39�F�!����!�������%�2L�6/������y��HJ�R!��	6��m=o;$T��_Q���3�������P����$[��K��	{���^�Nb���אk$C����"{�Dh�ˌ "�c�Jsv������"���?��Fh7�X�j����\3+f�mH�"5`:��G>�f9�x���:J��V/�S�7����A�:��z�X H��DSM^����k߈�q��VKn!�=�[=B��2��n�������Vk�&+8]7��E�j����u�@���}gL1����&�/,�חi�.�O�ɮkZ�E\tǕ�[����><�6>��n*����ދZ)@�b����*��Z��l��H�(��Q�K~�����}P���?�rj��I/&�B46���Qv�$Ew7
����e[>�WE	�pQF,�)9� k�u��rߣ$e����?V��rFͿ�SU��L���9�L���ծR��Ī8j˯�>νs4d����#}@K����9ڋ�Ì�0�m�{3w`5�c�ϱ�T������K�����8�+��ۈ%xe#�n�Nd���!a�Zj4^����=��NU���~w%>�f�.;�$���%-"9$�����U;����P�^J�M �$���&	]'����x��S��0����cˑ �I�A�a˞g��^[,_���F}k��x��QZ�G̾.z'��E�<
��y��oV�3�< ��|+�A��:syq��t���P�� diN�E�����	�f�F"�1 p�.]��@P0cy�
G�p�7 �|��5N�f���eIO�깛u��?��:U��rVr�Bim�����L��0�JF7�"0,���_��"ze����\���oH�b�e�8�2$��=��q�ۂ�Ss��u?~S?]������N�����~w�M|�?��p�}[������,_����Qk]2d�3R��ǲR��/fWj�/�����t���H'Z@bp������ї���>2�]�gDl��YDA4�1S��L���,��e�7�i
���O;Sa4^��s½�n�q��\�k]:d|�a�}NL��c�T}=e�����E[�D��~�� �/��ѽ�!�q#+�A5j�����0��)f̬�d��}�RܿMx��3����lpXvw��~V�CB@#�
Ѯ0�j�P�j�^�U����-�7�߮KZ�8ծ;�K�YV	�����_�@1��>�Ho��eI��e)̨��\0^��!~�dh���3c)�5�3��?IWh�dōAN� �!<��C]��ô�⻲- '\q��/���w6;3�_`�|�n��tU�Ic�;>� ���������[t_�#5}�F�KT��?.ᣉ{�(�	w�_2���H�~�G2
:��iI���-˪�� �Q�G�Enp 	���s͛0߄W�ꚇ�W���&�5���+v�{=	���>A|�c��I琸��P����w�]�&G��)(ʴ��y��	���tן�䚡��4��%�
}5�b;����L�r���t�xͲ�4"�|L�P�c�~�v�Do;}���Wg=���?��	�<\%��H���ބ�W�Aƽ�ɡХ��׉��<�7� 4KVM�8�'�IB"�p�O)y�w�)�G�P����~�P�%��ڷa�K\g�R���槆��N�IT��#�~�e$���Kv���V����v�\� t�X�<����!j��N����L����M�TQ�[Љ�a��udb�[m=�3 æ��`�u"�}	8����u�6�v����[�C�c�^���,N۱�c���g�����SU`��)��ؘgFՏ�t&�c�B�0Z��r��X�wnP�>鉞1��,U_��Zt�����6�E
E�Þ�q#$A5y��Bc�fO2���4l'�M�qW�M>Χh(B����H�ḿ����(8�$��
ZR��7 B���y��4ٙ|�$`yq��)mX<��S�����졢���-bD��_�
�q��t�-
1�<�2�>�J�_n���4�2�X�9%l��:1yъN��Z8)�=�kL�W(~������/R��Aj��lb�����G���T=0�['�����3ve{E��YI7,���n�2�JOv5�;F�gh[��R�
���B�|<Ϥ�d�3 j@+�d�U-��4b��.�1F�.1Qdt�4���|�-�e-d�Эi���t퓞;�w(�L"����U BxI���0��4��Q�4:ZM��d�dҠ�&O���G>���P;'hulr��� �e��B�ak��zP��뼜M�����/�#���F/�":�ɩ����f�n}��������[�=�k�Xl��I��'uGbb������M�@�u�����m.1e����}8�����}Q)�gs}*iȸ0���s������i����Ɣ���F�o,�2�4�9Lg�}K���|V�n����a\��f*#+:(!���_�0�q�?��P�'qEۓ�2�v�ԝ�3f���8��;<M��XN\�18C�~A�d��3>���tr$�"α�i�C��������=[	Ş9�N�M�[a������]`rXK����s��X��7�����m�zPk���r96)G)�:��E���1?�_�{�{!������%���:���N])��j������2,��=��� �6���4�F�9���|���s��"��?s�Y�M�41�X(�dc��k&�ٖ���}l��<�4�I�\Nc���f������`�Nߊ�;>��N��x�[��t���K��-�WqA�±CǣO]�\c�QpQ���q[)f������8j|�Ŭ���T�Z*�@��`r�S���t�is�!k2'�\{��ޣ�H�� 悿�����~��AM,����Ox�;�-;��5V�$�K=Vg�`�$:�FX{)�ϭ碗���r�;�&._<��VW�:r����FN��_?|�Fs�mp�wF؆�P��޲���M�A��	<�!F�r9�0�w�	`<�~�G���C�V�P�v��$5���tY�j����%_P����־&YqpsKurL�bl_6��د��1�n.�x3Q�,s<�2_锄7Wk�Ģ�5�z_��͍rL-�"[��a�j��ȓ!����� ����*P = ��z�*� �?0=f���E�l*kű�6w��h�>?�����{�^�¤i�� ;&չ�̌�/���P�0B,���v#`��c*t��X�)*�v7�6�;+�Wu�i�e�����@&k%Ľ�ó�eO�(l�E��?o��I��)<䩚�9KZ�o����[�����:�x�B{~+d�mg�ƒ���S�(�up��َ��^�~�B�V�+�����=Z��y��N%ԃ C��u��,��>�M5�) ���1ϱQ73�0�@`kk�J���c+B_�B9AO2~������� è����TC�k�P3��GJ�!Q{����#��Z�i㪈�֪�\}�Tgǝ�Z�� N�+L,r�U+:S��+�~'�N��~f�\rG��?�&�;f�źYo���]����o�G߈]��� ��8%Ӊu����Da���#�	N�e$J �}��6�J��U�d��C̤�Ɍf'���B�V�����G�ĭZj��*�x�Ru�e,]ޚb��F2��}h����`B_��1"��@��g[#�
/v�燃�w�sJ�>3��e$��>���2Nh��.�Pg��đ��[��m�V(;�Y)�]BO�)]>.�.�b���s��^xH�9D�ჅEp����e�{�	�N����p4'#1(�L�D4�Ib�����[B��2!4;�g\�a�!d�T�ȵ�6q$�O��]�l�(�tȦ�H2aO��tF���d��8P�R���J�d���C*���;j�(�]If�w�x�v��s�h%���D�DZ�����v3�h:�)Qp����3��9C�n�%o,v� �����K�\�"w��BI۪H��|}�P�Z�u����A������$�3f&��P ӌ�.���42Ѓ���Z0�w���*�H�v-��{/M�~"�*p]�Vϋ�C$�z�xZ�Ɗ�%&�*q�6)�8���PE�h��@�U/�p�b��k�Փ>.}dS�}p��ݎJ����7��'L{Ȉ}.����ebP�oF�Ip�w�^f"��;�=�v�o��'��0�&?�[,�C����v:N��2�a�t=���c`g'2:һ�d&�Y}�k��)��p2Ο�����w�Rkez%�����f��i^K�>�D~m4�`�1�[��
V�yN�	;�D�`W	�z�M���^uGlډ5%��m��`�-��|Z���/���B�}�[�1^g�t�1\2v�Q� ��-�I��"���^�*��;��/<�:e�I�cY��nLK��@��޲��Y1����z��q�I�z�h��i�}.p�ʴ���}^@k��z��̤�v6�p�������$�*3�������8!��6S8�\+t'ܔ$���3�/�e	����)Y#���K�ύ�--+� P�>�ױ%/?"6��c�C����0�1�%���bC�ݱ�&���HZM�����'��S1-�eP7��V<�~�� ��{?p�����֐����"n�^j�w��G�Up2�lY��ԑwg������������p�����3��E�G4{�$�ZX����(��Z�+Z�,`$kC 7��^�刼 6�*:�L�#��ނF�A!�ngU�{�?����71�:ʭ��c>W�Sj�N��{mm����LKj���FNX�(�8��o"���$7����y�%�j����!C�����%�f�ð"��1"|śq�ф��S*�r|l�`�U����;�k�.�b�dI	�%��q�c�eV�]⊨���)}�ѝc(�7 ^��{�q�+'��<P�K�q)���L��,LI�`|�0�0g�Ր���BZ#�&g�<B(IRA�u��d�7#��i)0��5�nqV5t8�FKa��w?oo�%6�e�0�Tߗ4����f�� 7���T��<��� K
h:ɰ�v���;љ❭1ޞ���@��u8K��j��ɱ���M$6����9p1ѿMNP��H�Q%���ߊ��A�R�Qw�9�9���&]�u@��f?���4�.W���3PFD���'GZ�k� �{��� u�J{��$�'�m`7,���N��B��h �M�N�O!���no9ߚ�j
��F����׏�;.9@o9����a
}a�E��:b	/s���$����l���^��̽�r�N�����s��~�@p趌���F������]\�3u��-�o���-� P�8��H�
�" �����i�˓g�>�`%B�v�wNh�P]�[��s���t�`@r�w�|� ��ׂ�o�5�!�D�0fmTz5V�����8>﬍2&��� �ۈ�*_�Qu*H�����a���.�p��#��H����`�5ɧ�{��҅rg^.���p������zH�f��R37Z\��O��ҭn�i;O�c�4��J�yǣ֓���0���}��>K�_��Ağ
T�8GI�_}�c���2�b���!��gkmuZw��m�J�wWQ)c���5��ԥ�҈�|:�L�ؙjqo�����3FgsXY颾��lR���?�G�X
����t�~Tո�!r~4�8�͉�dhq�/��lv�&6^��|�K�\��A�$�x0�Tu{��ܢK���~)"_9X �;�u�.I��MsW���T�;s�tM��T�i�����c���}��b�:�?a�@�����34{�������p�-���F�V�u΍��H^Y(��@�Od�EBG��Z�t6�_y�����(�H"^釨\3jU�&S�IzT"����X���'����/��J<=�}���`�lݹ&m=O۵���]��rpI�PG=�5�D��Ɔ��p�U�v$WR!e>�l���fEC&�� 懶��؝jF�r�s�6��'���nJп͐?B���Q�Z���,�`��~�1�zF4ߜ%n6���s�ypR(�ҩ���ߘ�8�����[��~�A��3&vdd���ؔ}S �D3��!��(w�|?V�>�������Qm�~���w���f�xvx�.���+INɋV�	�a�0�>����Ȧ�ǫ:���(0z�rca���W�0�T3�^�2�2�1Ph�^�;fj#�53~0å�c����Gި������ov�S7��x��	5=�d_Y��f{�X)�ܡ��*r��N/�gU�]�b�3s�]��+�|���Z��1qF�����T��xn��A�s3v ���@.���n�|�LW�pl�E��(�|�S�35,H�Fg��,����UJ�;bY�[��=k7q�56���P�\*ܲ���\Nꘟ#2]����Ep�bL3E���B�p�w7:��+�d/�!-0{���"�j+�J���^7�%2�e�$K%��Q�0��y엑�ڲW��/pO}Z�%`�LP������&����=G���"}X�t��r�ɀ8�
fEm���B�d���f�J?�*ܓ�d'�w�:o�m:R�3�Z��$a�|�}�|��!6\����+F�R�"�b(),S^A����M���(�}9�Ԅ����>y��[ԅ^c��H8E�}����@i0�ٌ���E���u���N�ZN�3i��VރP `;��Y��^�jH'۲����9|ٹ�ȯ��n�Ba���;gA(�w;&�b̪�DRd9���.J�	�l�÷=����x�����������buib�ZÛ}_R,�|H�z{2���D���R.��>�I�1n�(���>�R׀`k-�X� �X��|< x����$|��u�[�ٝ..�-8�ȃa����Q2�&�!�q��BZ�v���f�7y�#	�=(�l��p�l��xa6�rH������_ҁ$�1��Xv�^�>�J��1j|�m�'��������y������G�,<iKs�A�����3��~����a�1N��f�<t:E��z�vB��m�()}�� ��j}����P?�vXf�q�O�-�6.�F%yd���N�Y^��N�G
�Sw+���X��!_�S#��KP�4��hGh��5D��|��M	��?�n�����]2bs"!�@�x�'�1��v f�#)x�vt���h��<1Me�����"P.�q���}.r`a��ǡ�۽��(6~�M�G��˄��^[�]zg�|$g7؎:�[q�a��ە��%������'�����=Q���s�"�?����M�����h��	�O�g���w����퐖Bĕ��>�$~�g-�\�bWkM��Zbˑ�c����42,�T{���x`�2���L�ɉpצ)�ߒd�L/�>R]֯���@�����$�4-"}"|Z: �$M���_$�S_�4���;H�ƫ;t�h�Ňs�fj�R����~I�jWW�6�I��k� ��r�6�:Oز(&h�1*&u���49��+���I�{�Y�;�N��@�<M���"��"�X��G␄���WV�r1�2J��0وR�-LY��q�8�����ɍڙ�����@�!Gc-`��h@~A\��&�qP�]�j�bx QX�E��r~���*>#����"�d�<@�ם�<�*�"d!b+Fa��@�J�&�5�P.+���*{��0���NK��Z$�JYov.鐣�F��S�ϸ¾f�q2�ޞ�^�F�a�\4��_���
*����U��a�D��E�E��6�o��m��'a��1���N�9����h��NA1��ȥ�|ș�݀Aa�#�1PW��\��Z.�T� ^2dКkl���O������z�/KR�������D��-+�b�÷�vY^�[�w?��G�[yX���j��N������>
~��@!֏sJ���f�������6,|�@��#BY����]!!�Kb'�Vfk�9b',�"j)lΜEu\�W�ň"6�ě�����FY�w�cmg�A�.�b��~�a�5RP��F��3�̍�>�Y���4��ҡ���~j���>���e~8��"C��_��A�='�=���6��m�shGQ�}�w���w��:n�ͦ���(rɀ�fJ��i
'�LB�i��ݹ�YH&'�hNi��<G��\�@le&�Ƙ���&��j�w�mw��l��`a�Vc-I�#�ئ�b$��١�9V� �ә㈩(t$|��F�*_���)q��{�������W
�k�(l�T�)E�\Lq�5ř��j�n[0U�'t�l�Ç��E\4e�$,��~�};z ��f���aƽ)߷z�⹤%��2��L�j�[B����(�[j�@��~����u���r=�n���Eߔ�Pm3A����+�폟�i?����r���̬��$���VC�x��h4�2�^���/#��4*è�)9��n�	����kp8���.f}�6؛�A����s����^������o�[��D�O֍(�,�H�����J�����{�&@w�+���>?���t���&���@n%F��d�Կ,6��
�	⤾���*-�������|�9Fp?~x�H	"ڸ�Xβ��>V�Y��6��CQ?IR�r�rX�6 ]	�鮆�����֮�U�17]_z�	�-os�#�g��h�Ĵ���yHD�\	�Gn���Zm��� +w�sXw�O��z6jJ�.g0)w��-�Dߏ=��M��)�r�48��*�D+�h��J�R���}���O�"��q��yl��"ĝ���}�v��b6� _f�GT1�~�E��}����t=����O�= Ĭ}�����}M;t����G;�^h�Ę�4�ʺ/i}!<�s ����\BӋ�-��R����0^��S�	�V��l#I`n7����D��ǠYU��gO�Y[	`Dmx�F[��*eARa�]�/�<�sƛ�c�ل_�arVK͜�5�[M	4~�ѱM�{��3#Y7�UF`�4�,]�`� @"Li���BС���Qt��d�O��8��C ��ݽG�Z�3��{���;�U��>���e�LENv?����#�x��D��w:�f�|���L�co�DYk���#���L�%����-*�������@^��Ց�TXO��߁��1$E�E�(G�[��/9���n�l�i�Q���14��nz����M����̼��f�z�M9����)�G���np��gt}�Ϊ�Q�����gC�p��]����X�/��l4%~��O���3P�z�}~�P������ �K��w�F���hG�x=IX�.�@9���y)�o��Ir��Q4�K?�y�ɝ
+2��'�7N����ռ�|�;�]`7��V������6!������b�8!�,�FEX�6���U#מ����VM_]p��ҡL*ӷ��҃hQ'ʷ��a�s�_)-
�r0-��LT/�B�shѽ��cO�A�?;c����bFJ�ɢ-�?|�L�\K߫r�%��f��%
Z��w���a��`�ۘ������A���i
\T��C���8�3�X��`0�[&�<����v�vWpD��3��$�?��J�_!^~��$�Z~�0|J:��=��D�k �v Bމ��� 4b�/ϓ�$Eۑ6�ykI��]�[Ϫ���5��os����]-z�����H�8
���i��W2^J=~��V!�u{w���w"��z�.��p��L/A`��e��$	@!	!� �6��@T0
�(){.��&x �T�=���~!e��S4�s-���a�*.�,ܰ���V���H�*�c4@�5�蜜}�>��������_FEKQ&����r�I�����|��;)�����y�ĵ`]e�>@>yS��O�>���|���#F�㮖��+��+�F3�����\�<�����ڨ.���X# �m�S_��m&qD����V�^Z<���p���w	����d��v��l3��/5�|° �X���p2n���a�GKGM�w��'��2|�3$mE<-�k~���C�1����?-�={i��R���Sj�V���yq���]N�v8�р� E����l�l��,�~r�A�v�x�h��Os�kI8q7Y�b&� �BR��s!B"���@)�惗�������uf�Y���ͰMb������ef_�>Q�� ��Z�jb-W�&�8xɎ"�B��;���0!\
{��z!Z=�bD�7�[(P���7 533(ْ��N&^1/�Ů%��/c���{�S�O��~�Q�v s�˪�}��d}��<���"��K�z4,3�Z��J��L��n48���g�)����w�����C"�'���l������
%[!M����=�/eĶ�����梼�O�y7�D�2�1��[��. M��ޫ�:J�&*\��gf��V;C��>�X&�<4�3� �㨘���̦S'FO}w�_6V���
w�G	[~x���Qu�υ �� S���W��>{�5ڻK�I�ޏ�U	k��C�AM�1\߬�|��d�ދ��d��-��p���i;�C����x��*���s���-΁�WY�0o(N�l5��V��I�=l�_�1z��t�2}��5;n���L<���j�Ѳ�A&@&���*[�d![9�k�9v�T:�a�g���S9�b�e��aO��8��)D"���ඬH`�������;�nt���E�@=P�YsZl��~�]�)G�.SO�����Z������Lia(OK�{�=w-R����ǣ���Y����1�� ���|� *�XW�<$��H���U���h�4 =���+/p���?���9x?�h�Y؏���y���Ho�B�%�-�$O-g"N�&�����d{�n>4b���`ѳ��*RI�}��R�`�r�M���e�J���Nǈ��!�r���s����PG���v)����m]��-N?�OW�����7��O�I3q� ��m6e�`� ��-����o"�1�h���q�E2��t���4QUx牋��3�u�^�0��^0?Fd�O���!Q��I�[���i���s�袦T�;���ʴf��ܜ��[��T�$�V=+����5=t@$��z
���������m1�RZ��������g+9��d-�̐�b�h:�}�ɭ�R6JkQ�����[�U�Vr>a\�|B�4�#����TsO���ßݳZ�DG{����*#��
]�Ѯ�o)#�)~�J��_� ���"�'W0�J��z��c����'�W�1B����ޞ9H{�!E����oMC��F1��҄�>������B(\��2�Y�m|��1�q�vK�=��W����zR;��j����O�>�/�۝��Q�1��}E�Fk�������N�8Foj?������~��瑘8����r��}R!z{�<?��WU��CT�h
�ֱ6۫���×؞�?��J�0G�
H����ư�zK{�W�7�j�j��Wå;yD�A���͝�	�t:.�kgΠ����?��歕L�N��Ri������ھ?T߄� {2e�]6z�3�G�w@�!^������[3����댵�I��'��4${k�q��R�u����U�A�Eۼ�@Q��i 	�G[�+5�V�|=S!�Oaf�[b�$_�@LkhO�pU!H��Gu~�pƲYet�z��tʜl}L%�����F&����<������5���@e��{����UP�E��>��\Ǘu$���U|�'O>��:�E��M�t�*��Fʒܳ �9m�`��
�cS1tJN��T�p��$ ����yxҕ��Ў��}��'�b��w��2��,�f�� o����|�{A�.�pm��`<�U�����Q������(�*�h!A��6sǸ)�Q�~O�3�9
�;غ9T;���k��ɆR�f;=�ru�;^�Ϊ�~���
��`��������6��Q�@�mW�px���[���2�8�UE��]�����U9ی��'w(��W�1�Ҍᥚi�R��ܯ4e�|���]Nc��c����3|�y�������A�n�8o�a٩�-a��~����~�&e�l螳�z���X�W���>�����'.-ִ^l�`��S,I8�}�&�>�+�k������?����4���3�t��n�����a/���7�\�O��,�eJ���ᚭ��Wn��v_���0ys�sEӟS�73�;O�aZ6qM�gTvY�H{��(oٞ��s����'����ðN9B�J�רFĢY���l$�$t��O�zuY�n)�1V����|�����I������`��p:�3�z�����[ȋ�^�B%	�:�i^i<D�%�͔��\���79�aKW`����o��%4u�ӦG,�ƈk�O�ʈ��iv��$jI��Q�p�^5Q�_u8�@)Gba���$�H"YJ}P��Ka�D�}���Z:r��H�L�p�u���Ѿ;Fp�gax�����P���iD
~a���(ϭT#
�1H�.�����EǄ�#��dӊ����d[��8�?�jq�l�1�S~�(B~I�6�A�)�~J��$�[�f��Owc�!��ڦ�Ña@k��;�u�b-%�'W���j�jtc1��Ŭ�{PR�̝��I��E&��F���_�B%��}>_Z/�cS����oZ��M�T#� .lL(�ܠ�M_�o���������`�Fl6�a�bs�2A�kd@�E �楸ӧ�����o�������!i�opi�*stWN�?��p05qK�)���b,p�,S����!�q:����l�V7����� 8:}
�OBn-�?�5��>�Q�&��O֜ؒ�C����1�JɏY��3��|&�wȹ���5$|�s��6�1 뚚�о�ONˋ����ԓ��IU�`�mI��~gH_Q���]��ϙ\*��׌
<�o$�ö�Z=1kq�j�g>)�sb��B�:z|�"4$s���cO�ܣ���9~�f.�_��� ���H��*��oQ Ӊ�I�d���E���l���t��M$ АZ�`���l�����1�`�(-{t�GT>[3p|��.��7���tz��t�v�p�}r����E,����B�t��)0!�8�%�~(O���2�*��H�Y�D|������l�U�Ѭ�Q�s��k�@��spq�u�X�I�>
hu�疤Ue ��q�[x�*3��.��K����q��?��2��L����]�G��	 �%0�Ա�>��4�R���T4փ菶��V%\I�Mh��	h�8V����H\)h2?�DY[W��F��Z�I\�)R�Lά�ˋL�Ir�3��ʫ��Dy�=ZY㓟� �����cxR�jP�)8Y�Շ����ǚηG�m!<r,C+F;��|���&�2���
?�� K�t�#6�
"U����Av����k;��(n�U��{g��5*M�6KlkS�;S�}g� ����bm]�XF�!�o�p��/&�hՒZ��NX��6��,��{g�UZZ|s���8����3ͳ��F2�a$�kW����+9�G�>��'� �\T���qQl`�.�N�T:�H��7݈4�G~��$��^�����f�Ƈ���|�Qj&��bH��|�Ri
tj��i���B�D�aV���=�zu�x*�۪'Ɓ�?�ؿ�_�7�ɄK[��Iqs9�l_�ei,3Ǿ�����뙌)�m�5��ɶ/�����X5�c��Х��׳@5��Óe{q�]�O���)��G��־ca���Y�d*g
���g���~g�� �6d9��<W�
�x��Z13����М:��t���\o:%a�|�$�/�h���rq_���+;��,������z�PI^Z�7u1�~�&g`#��dDd�l��ɲ���:$:K�Į��n�:���G��Y 4w;�0Ήo�N�6r���F�1�a��\����EB�Y�>�-�M�O'+��n�6�p�������_�x%0\1^�Z��0�]Qth�T���j��[�P�؆LX%*$�y�vܰ�U�P�
���K���ZCN��v����n���L�1���焞�����pY�w��9��j��=�;�0He#~fr\c4CΑ�A�p�%�>I���BX�OX�7���o��̎���OaQ��,��I*VK�}����֍=��lF}?����h9��X�^�޺�ݑ.'05�I+��|f�u�G�"�0x�������k�e��DE���k����,�F�jO��f��P0��ܾn�RQ2�9�5���-{�;^^�gb�嗠�d]D���������;��m)V��V6I����Å|�/	ŷ9x��-��Ƹ�O`��>����u�~[�����ێl����U��Â;=��;�͑m5(1��B�1�
��.��x�h�~�������t�i���&��!�r��)!�:����׭���,�p?�[$+t`��[Fm�!�0�A��q@j���+E���m�tȳ4���^�1��$�-$�Ett�����a�Մ2�ה��a�u+�� KsP����R��FX�PK�+�ǩWf����7q8*���9t�Hr��it�����pN���w;����iv9Q��.he8 ��b'��X��2�;T&19��BZ�zod�BFT���*���ュ��m�Tp�ל(��5�L����f�%'4��h|Q�/�6��t/���/@�y(�*Mu���D_��l��GKy��=Fm���i��V��e9��k�B��λ���	Yq����o�cW_���� ��aJOlk�y���m����&#�U�-��<^��i�V��w��v��X���}ǫ��IR�Yk~w�CM�Is'�]��#혨
�^ħ�Ew�����K�²W
ZQ-���h-��h��ޟP��<ac~�s��;��8��f0Ўn^���T������1X�<�s5w8���vHT7���^�C������HJ���gg��?9��0��W��V8v���S*�i�O��,.7I��Y>>��)�^��}v�����r^���'i��{��~�sz#�O��?�*/(�1�#cr���f[c�ĔL�2�����`V�i_CcC��P=H#=H%����.��VÃ�'.�9�����J����l>vp��auq�gP �$�nѦ:�ප'���-���]í�Ɲ��:��ㄣ�d�ieR��j�Z�f���
44�����;���d�Z�1>����ۖ/���7�
o�:\�B��/�����s�|�����k�F⹼q�@�6�ڻ��If�lf�g��3Q��F��yF��=���?k ����ޙt8�f5�и���]]q����h�E4X��|%ѐsIN�3V'\L�zƩ�.�+������|�̢"W×�/��t H��J��\1z$y�Y���qD8�LL��&L�;|$���yNH���1�J�R��X�}�����6m��ze��5����bk���}�\��"zUM?�=N�,2�G��ҵ�dޡK�L����
m8YR�z]���U�U�g!�(��.U;�����
×���ot���s^}+ k�>Pf�i�[�Z����7�6�����I%���up0�t)�2C2�V$�.	K�< �`9w��-��|0w�^��̓��2U�l�X�_Uo��	K���	
���,q�2C۶�R��M��/��]�!��]S�����|�\Xb�R\E�,�B��s�����i� n�S��Mq1����y[���9؝�7�ZM��A�8���ܛ��� �,"��[��ᐪf[˖���{�{_��飏o*��@�Ҟ�I��X��|��t;��p�P��cK��}��=��B+TR�ȕ��Ӫ
n� l/�� M�5σ�:j�X� pp{����uO�A^���)8p	�������.SD���v윑#��u���͡� y�p#���_�q�'�~��u>��O�=�D_�\vM]Uw����5n'ͳm��q$dGA�I�����ZU���0E�܌�YP=̗��UG.zB��!>�c��úf;̓F���8"���V����k(�����<;�4�Ѥ��(PC�����B�#�Sz�#D�x�a���O�sP����䊭�4�X��!�]��Ī�xzqv��^�p�,���hf��T�]%P-p������	5�0C�:5�&M�K����OC��n�a�F���0ޢZ��Dz�)� ���wR`�c%�;��q�7����*N�QPB<b�d*�j_��V���E%^EC�[q���w��D��7����4��%�����8b�|R�nW�U��5��(������z�-g���M�k��U+�d4
Dn��a�%|�dԣ����\~1qE����d�Nα�uɢn�A#V�x1��X8��W�VZکg�����Տhզ���S&g$���5�kH��KV��vh1��\�(6L��/�C;���ֿ�;������<�#����(I��I���z�h�V-bI�UB��"��ϰ9�7�)�� ^��	����`j˃�D��.=�j��?�(3 �����d1ҏ��;�/Uď��]����~bI�+���|�ٓ���}_K��� A��{�;�lg�ʎ�W���ċ�S���Y ��&r�MP!X\I�q�N��a�ן5W�dN�66�D:z����tJ鬴h�+���^y>��"�KT�	�9Ɯ��4JV-���kO���]M���ư�$rIw��kѾ|��3s��h������%ߪA<t$�#'�̪y)zq�Ѳ�n�j
h%�[b9��n���#4�4��FEs`�,uˊZ�Br���u剏�q.�7��U�%�J�5,�:���ߑ�^_"Wb�/�7�����EQ��M;:b�(Ȅ�DJ	�P�qh!��J0�k}E$L:>E�/�n�^C��Q��X���U�j�xt̃����RX��#.�F��`���j�]����Up�+j暉��"�_��_�u*��w���u=X�&ENEe�/��g6���x�G�B�<-�h�|�Dj$�8��݄x���y�R��}B�߉o��6��i�X�9�`��E�<��'���2u��1��۶�l½�X�X�.�P��=+�9&{�ܠG9��"l�ZÐ�h�C~)�-^)�������� �����i��.9�k�� ,s0����,�U'E�������?9�.s>i_f#×x��Vwv~þ�p�Ъ\��0���o��')-��%�x���"iw�B�n�SWGp�f�(�UTf�K���&V�U��am(�+x!{HFȄ��|$ �0��H��V��v@���|��S�Ϭ	�Éh�i�*�w0�68������H[��zOJ�͙���EM|h���C�+�����1���~�~ǉc�?��r�q����'6mQ����Խߘp]S��?vB���n���՗�7�x���ٮ��v��1ۿ�ÛÀ���0
�������E�s������Q��)��1�۹�HO��%�Wz��ؕ~�i"�;W�D{�X��r�ԫ�ˊd����� ��=^�v��(��|k>!��(9��fքn�An������<�9�@`�#�Y?�z��JDޣݿt
߮Rw�<7q���S�m�K�{�:Fˣ\��֠��T�j�o�D�]�3P������������ahc�?�<��䘬1�7�gHZ����rg�h�d�"����)Ӟ`�8I��;T���;�Z�(вђ��}#eS����tq̕�3�	毠�)sl99D)�ZZ�o��*��H���TH#(���z|�C���	�����n_f3Vmg�mk���h�Ѕ�5��@�Cޡ'NV��4O*稷�c�0��j��K��֪����cf����8VA���W4Fq�Œ0��סN��M��O��xT���=(��j4�%�����;�l�X?����7sk��2_��q��EjV���<9�E+�K���>B�����w+�St�@�����2*�a�����l68Xc�dL�-��@K��� �C\��_�>��N&�P�Q�t&��+��e�e��"_6��FI��P��A�nhJ�(����4�:��DX1_�ĩ5���G!]3�`�!� �fzZ�,�H{�¶�H<S��2"���붰�w&�"�7��	�V�."Ø���i�f�A�$�Qm`�fꀍ��(�A�B����;V�?V��t[��4�2/��^HM� kYhC�L���|Sq^�����*��zʶD���a�~񓪟��d���aUWG�c�mp�.��^0�T�V`���d9�I��	��f:���@7�݈����t�O�wO׬j���Јߑ12�����3|0�M�����p:7�K��VT{uB��u6?D�k"�Dw﫡����UX�ŷB�[�^u -���((�@Rf���p)d���J�Ѹ@���
6^P𱨄�;;^�v����^3c�O> j�q�7s�Ջ�����a<�P4֎�[sN��1ϱ�{�rs�?O|���{�	 �w��H�`�k�������Y`
6f��3�*�=��#QtZ1��a0c��M�!���y�s^�Q`^Y����DuI��'y��mȭ��|J���_�}��ۗn�b���򱰿�	L��>�\��E��L�����Y!i5���6�"��??�M����FCdH�}C�������Y�v�]Ær��m��2 }\x�h_��ۗ�Ts�����/6��g�ʖR����
��2���J�q�\Na�u�add�BQ.:��d�3X��ȇ��K�u������-�9q��;�D$ ���P�I���_�n���zk������> P%����K�3�a}��@�A�4dv�M�D�k�����loU��8��D���%�l��t�����,�T�u�_�^u�ҡ,�O��ͼB��������XyJlS�N��d�׎��C"��p�o7���u����I���t��(cb��ʸ��D���n�7w�s rpY�@��*�Im�R=0ȱ
���|fԢ�S�Ԑt�����d�w�%�7�W�0�l�{)S�9K���A�z��zrD/��񘌁��/�m:���'��#�H�����>�w���^�\�La����u���pgb��=��5�@;n��� ~�1�z�aM<r������Bs�����������q�_J>\��z���>=Js&Tɘ:J�;!��B�B���$�u ������}�|Ί��F/�s�����Ϲ%y����7����5xB�fo����V�ʙJ���e�&��ב�뢲��cĎ�づ�[J:LGgg=�=���^^5�k�*<Ez?#�&"tE���С�}�Uup`�vIU&y��Rș�o��Z�+��U��.Gd;�V�߼fS�������n��X+�~���矔�H��+7Cר�\J6g+Ob1�OMK�a�˧�A���՝W��f���F���3�!��H��7�."� _��Z�c��b��s/�kV��#_��z�`d4ч����u-�P�h|������c�Q���)��E��?vQ�(���o�P$��@�ҴO[��}-3O�S�@C����� � |7V:(���ݙ�̚���6*�26s�0�xyMx��ޣ�����咦��g�Ր�G�"�$"G1Hc��2�O[b�ϩ�A�ĊJKoC�9xjou���ܫ� T 5��	L������������8�5�2z�v��_8R�Ǳ`/�͝���f�"]B�|H>��V� 3:"u�X&�J'Ǉͭ�c�V`��^�K�C�A�;M����ͭ6��NF]/�U�*����h�xHX\}��/�����Q��n�ŷ�Ng�!��$%�*n���[e4\�R����C@3�פ�S��.i]�A��QyZ��%"��P%����[��](+�\�<���#k�S�xƠ��@�S�3���xUөz�K[8"�R�������jRü�ެ�:�h�_���	�r����ODk�>yg���޻��Pݣ~7�u\b��A�mJ.�KCz3�K1�}z����ӎ߸햹�őCb�J*������G�L�Z�}��װo�e���_��������&��A3*�*&$&f,X���ϱg��<�}����)���`�:]��K��rJ��\��$�r�_ J��?I�xi��#�F�3*ܕY2��.�j�J}c#p�m��ԙ�d���O��V�\2��v�}�[9�f��)�A�P���Xk�����fn6/�89pv,�<�/\U}of>{>��I���'u3�X�G�}|a��Y 
�8,�m�q�hl��5_*���YLܦ�Ch�$>*�������s�Gm��!]C����U�Hkxq
��y�A�L0��"�Dt�I�i�U�~Y���iu��f�J.K�E��y�����PU�$_z2�z�D/"��������0���U���o`�0W���q]8��~ ��Y�o-�2L�{�w�~(��"ȅ���VȦ��])����������~�x�sj*�}��1'�Y
>=��z�k�j�q�A;�R�#�$�f[�h�Ztn2:��BB�5��M�Vc����_Dwy�(������v0���\a$u�6v�aL����0�ޔqQ\%�mݍ*3��EҝD5],��y�o�����W�2T?:7�%d��p7W}BD�>\+wd{������I��U���Z���qzkɡa��c�P�}�oa��I�/�-��Բ�9�m���'(�\�������萭xP�kn��#�����OU�41`Qƶ�fRЄN�WXf�n����;����G82�����S�T�� |"�bb�R��3fr�[�&����3a�(M3��3c�`(uO^
���~�	��)�
�E��Fa�z?v$���������i[YQ+'�l�Y����頪�h'���1�8�&t�1Y�؊��|�[���na�Qê.�;ԋoA���Uݑ�#UJ3�?��ts��u��o�1����(��m�@Pߚ�^���\S�W;ɘ��6/��Gi���gup���\s�ߺ���c���j�D����2\��4U����"��-� ҩ0���%�iRFٱ!&s�V�T�����KPĺz��^�*�z�e���K��K�J ��� �Y�Bm�~�ti�ߚ��!v$�x9�w�����Al��(�Z���Q��f�=a���͜,p�ʫj'��+��6]�2���
�1�O6���z}G�(ef�N9��VM��t��JS�3.�����N������#mV�Y��Г�WU���Hn���o���t�Z� �(͎�h��/��p.�k��G�kf�cѴ:��Le]>&
0'^`��ٵ����t� !���ud��H{2D��8��ƌ5n��G������@�W�w.-�	��HϤktܖm�E:�5f_=�jWZ2�<e��'
^L
��yn�[�n��>���B:��5>1?�tXn�1͟al�	Ŝ�B~���&�/���F3�����$���&D�WX�5t@�ޞ#"��j�X�>�ހ3�b�O�ws�zCa��_i;�'� 2+�LͳŢ�??�f�����z�n$�Զ�+����Vb_��z\f{�$�ٔA(���9v�=r���B���$E� ����9g�#��h�O6l���?�`V�^�aI��n�0�ۉ˸v��l�7���wć��$dm�雤s%�O�#\�҂:�1�O��x�n����c���{��XC%���Z�����~�)O����h��������h E���K�v��^f>�V`
�o忑�Eʏ��&|�cwb�i��s���DF�o�f0�h�n*�;.a$V�a|�fb�%�0++���d��YV��R%�K3)��m{���	�������q�$)��ٺ���
�.R�D1�*
�`��iH�Ͼm�n��	Jh������Z�΢3��r椏I(L���8