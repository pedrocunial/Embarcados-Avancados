��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c�F�%������ !t����<n<����3�4�VN��@���82e���y�N��!�"=��/(`D3��L���|�e�S��HV��&���Mz�A�F�:;���2�Ô`E�֭>��F�)��&0f
�n�q�f���G�W0.����3_R�\�����J�2Y'��W��ݢIm�cC�e������Ǒ��
 ��g�'ɪ,�x52|}�@%6�#�ɯ�n]K�fSC�Ǉ3�F.6.B�iKoJ��2��<�qVP���P�'<��`�臼��tkW��2M�X��c7�q!�_��_7��	������w�\��K����zlmș0a�m��Z�U��}%]��f��+�_6�6bb.m0<5���&�xǭC�GǪk�M��ٕun6㿜s?[>�]$1��hzog�R��"�nk"0q4���h���1��
*==����M[,��q��wm��`�Ǆ' Zl� �g���֬V�G)G���^��FZm�,L�8R4�2�긦���X�k�d�ejO����F��� o����͍��|�{�Rnk�~�=c��g!!���l���z��I�:�9�q��_j&]S%��1�CXD	bXl����(�'��Ealuy"ȅQ���j��lg�������C��/�U�9�"�ئ2��c�Ƀ��X�ʧ����Xg�2Y���/°;�u��y��&[�����[9FSqJ��*PyE	��FJg8x� ��5�Qx�Wj:6�`�j_��e7�A(�Z6�~�A> �V� �R������j����W0��pV ��)[��LꛒsJ�G�]ލ�hف����}���z�AL�R) z$N.Z�����ք�� 8�*s���	���f[�2�
yX�+�:;��یh���b��8�ۮ(6dvD��v��D#�-E����0��"�}��z�5#������0ז�5zU����8��S�e��=;oދ-!<�m��ْ�<�P�N��y�T{Y�`16#�O7��Ď��6{��*R��F��dP�;����^I��/Q��V���{�l/mG���隗֙^5���'W����r%��/HĬw����kw	�2�|�V��?%�&�Y�x��3@�[b�JkU���}��%�	uL�f8y�Qy�6���}��B�f�6J����-����ٹ]xy��y�>��N]�U'�����U+O07񷈷��b����7�	��\�c[�2��;��-�Akb2-|d�z:m��u���+� �+}}ų6��D������6@�e��"!�N��Fyn�;��˶�4�}����?�OS���ח�n����V��}{�u�$��YSZ�Y�`������q��\^[����u�9)�������Y':}"���xf��Y�	D4:U�#͹�h�c!�=4��.j��.��X���yy�ʢ
��O�X8�XW!h�t	�����lˋ�3��m��3���ߥ�rr�P����-�
='J�5�����&�"�zuM3���C�4�*M�����cu��7����c&��'.�S��;[�TQE�}��1��'�6�m4v�J[�T�d�� �E�X�E�1������V� 95����-#4�����l%��V������n��i�hR��֝'.W-ۂ��>�n+�^[�dF�o���ąj"9�u5,0��<`b@ܟ՟�	��!(c�v�,���x���@���l�yq�.��D�F�^���"��H-���(��ǺR�o��;�B�x���n��UF7�"��_��W�ț���X���~�Z�a�XPƴ�)˚{�����^���s��'�����g�=�-[q�[�������:������U�/�EK �fć���Ey�y�M,�K���,��[��QUc�wQzv�����dr�
��~��K��ru��Ί@_����pN�}���#����*K�qm�H>\f�腯��jF`�M�(��_i��������BSଠ�iFiOw��$��,������̱�-�,�4�4p-����(�W�U����h�N,�rУ'n�MF٦�\N�S3�D�b���#'��
~�D�7|��&���׸�D���T2�Z*�\w���?�mKj��o�gek�Gד|g���Y�ґ!H���`\Z�R= I1����ұ�`��kGFk�(�3��{�g"���e&��VY-�����kh��ל`�v>�t*�ݣ�Ϸq�+_�ܲÏf�#���h��BflK�Ѝ��RR��v��xi�g�M���<��*�}w�����Ű��c y���M���:y)�H����>��/l]-F&/��턒F{ݟU\9� ���1����) �4 bV`��̣�����×'�@5&Ν<�P�//�Ec.�:�s�)��������ij���8�� Ĭ�ں�O������.�0��>�����*��ܸ�4iu�Z�0. A\򘁺�缵&�f��S$쫣����l�P��zzWع�/c����'Ua��,�G�ܶ�I3\�C����.����z[�3M>[[:'/��j�����/�\w�����%^�FE.P@,�v叾=,�p�͏�����^��h�?�l�{,K¨{2�(���v������H����΀��E����@#�*#@�b?�p�J�byA�_$�_Lެ��3}�x�_1�3�`�a4�K��8v��3�|�it��Q*��Vp�[l�s?70�Ǚ2$#M~~0_�~XJ}w��ss�;"v]��N:�#��#l���q]x�}��
� p,�xUy���~��<݁�2
�e�/�vŜ�N>�H��UpO��{��Tz$���(���u3�"~�����0+�9��1���A�e2��n���o�k&P��Q�4�.
V�}�2�<���N��lϦ���yp��֦��}��5���e:{�����s��㓱D��7�&��0k����@$r`?����P>�A�K^m���`�J���y�B&�s~KN?���_d5��OS&(q �����GS;C_*YJB��;�
��?ԡZ�u�?�o�1��`z|�q�/n�AGk2:a�H��x6ႇS8���M2�����%)Jò[�Ѩ�����"�Y�� Az1��1�X� s��[�)|�US_�����K>d���k�r�`��8��3V��x'}&˝�E`���u���Tŵ�MԜ���)Y�Phf7�H�M��ؖ�%��G�-��a	t��u��6�JF���H�%*��LE	��p	sW�/iT����������݇?�C��f�e��g����B�2�����ݼ�������̪4��ְC˖��d&�w�^��ɠx��f~9*��[?�E`�e�8L&��U5����҂��چD (�U����D�B�x��6^:䭤�B��U��p`���!����y�lI��jD7��@-���İ�2(�Giئ !�O���4��c`{}>6r��{=�~���[��XqN��٬��X�/�@}Z;� V	$<����HA�(�RJL���S[y�B~X�W�A�Ҏ������5L����mKH�:�F��}�m��ܣ���~_�O�eV౎���²K�n��$`�{bd!S��|reD�v33���n�`P�d�-Mbh��\�[Z�'����X	I���^��prjP���ZI�|j+���x�" �����cs�����o���@�N�1�~iFA�l:u���4S�ڧ���k��]���V&�k�
l����3�� q�O�AXP����kE�TvA�?R��m��b߳u����~���m`�ʄ�1�Γ�5���]!���^��V�	��ӫ�r��@�T��$䮘1?'�nk���ɕȋ����;�^�*,�Y�|�0�I���1*�m�_�i�n�1�"�9��LԿ�H���=�,%ٖxɨ����d�~��W���*�,�2��aڜ�o�Ւd�f��x�]�rAd_!0L�j|I��k��.#���E���0Qӫ�,��]J�R]�U��y��FD���u'�����OA��õ~���͔r�U}�goj$Ga.3c��5Q v�(�Z
��|�N7����z�E�����[S�RN�%:w�gM����؂+��Nٰ��򪍯Q���^��SV�/E	�SL?�� �^u`����Hu2�P��4�����d	���[����t75����ѫ#O��@�ޅ�myg�U�m�q��np0Je�Ey�崯���R��4���=���0�BCs��A�$_��k$��RX�>4Z8E#����O?�c�0E{����U~ڞ)$x![ꇚ��O��)��=��j�N��[�>3�`�U���S
b�|�-�#��C��E�x��T:���6��~��W�1��1�j	z,H^��ut<�0Ƭ��#�=;�r^�Q����dm1���Bt7�����QŔW��\�dR�W�(o_#�E*Aڭ�:?+X���m�p�s�ђ*�m�š��lIR��B2Pc�'0�{"8����t:���u��F�r� �{9ù�N��)>f��/t��\nX�*�)�PN4zM\�����ɏ:�{�D�"t�<Q�����~�p�nΏ��C�2MWK�:�M�M:ђnҹ��2�+a�nl=��$�v��o��f w���
��V�9:����v�|���pHiX�|�\~�1xS�㾵�X�Ƥ�E�]�&���c�{|��DE�f��o�d���׊�g�uWjq�<�Da�(�]E&�~E�qB�y�Z�;�R=nd
�{09w�^��#ٻ��k����++sE���=���"�[z>6� ;��M4��у?d�^1t P{�-�p��י��x%
]߭|?����n����6�,@��:*N�Ě�G/���]E��xJ5�-_�.�����H_�Ȱ ɒ�!�ڨ����_C
�*+�Q�����n�:��W�S3x|\�gU�|~Ǫ��|�$���EH��G���U���Y��V�?(9��<&�V>/���}�0 �QDF
�_��Ao/���!��;Ѭ�(��Wc���h��A�d�Ӵ�じ!��:�|�F�y�:B�П��A!������*�[�0���牴�=��?xV)�e�jJ�m�.�c(�&oOM+^��YWL`ci[�!�*���A��s&a|����׻���F�(�C[���mGh�E�w׸ ��+�ji���+э<0�|�����mӭ�.^15@o`���%���yh��?XF+csУe���(��<��ö� �R����l�ՕH����tx9T��g��r�D:?��U��b��9M��r0��m��O���!8J_m�YX޽'��/`�n��6�,� �q$����fNܾ(f�1��G�]o=�Z����0� Q�}rɹH�k7A�a�P�����&i���EކpC���J����t��m�bf;}�Y������/lo�6�Ăf��j�xp��|������/�ǻ>�/d�����g$����)~��B*����,.@�Q�nR+��WF����7t�Q�ͯG!؅B�
�
��^O�����w������e����~t+�^�*^BQ��Mɼ�~*����w�\:�.j4>���jD;A���S��r-�H<.͠5��DD~le�%IZ�W��{�I��ǢRM,M̲����MyF
��4��9��S�* �Ӹ&�egQ1���y�d��%���y�>��u_.��,��y,\AV����F�rO�^^'q���}�Jĺ��|5�+�Y[׊�R�KI�=�f{�֖;T7�����w�Z�tK��~�6.� �U�q�=�3P�l��&��� Y��S��Wx���Į���R�����m\"�,[��.�E�?C�}�M4�,�*�h���PQx����APc��C2ɒ�o��g�P��'�U�Ȭ�`u�(�+�H�a�%x��s,7�Ϝ���YO�Vn��Y!�c�e��j�J�)j����׷j1u(��6AJ�x�5�?Bsﴏ��<#�	�]��WO�,���lxD���:�.3<=M���Q��4K�g�bn|����m�I�Bk��Y�ȑю���u"�z}��$޸����30��
������!�&S�-:�@C���{�+�4۠X�j)�e��$��,���`vF3y��x��,��AS���#���6L�`���]��΃+�PvClC�U-i�E��în�X;wƹ���oWQږ j�"e��g ���V��yև+��Q�u�U�~�"A
��l\�:�@ �U�Ⱦ�F�WP!b<���\���F�Y	�9r}�2V���.���]��&i\��hy�;5O���7�>����1�xD�:0���C
Y]R|��k��'z�H~%j0@G�=��׭���㹋�:*N|�����8�r��˞OՈ�f#QN�df��H.�k��Jd���&V~s�4oiX6�>��,`�k��#��T�j���1���F)����sHx\�?૏�/��IK���P!VH� �k�%�0 !x���M��C�Uva�а��#Cg�V:V��L�O�}��w*wq?����a ��ɿ���n9-i�Bf&(l�d^ɷb�!_Q)@@�"ZC�ÅX��V���V1j�3W����Z&A�_ӈ�`:��I
��t�q"�����X�_+	�=������}����:>����>�a5��9��6f�>/��>�v�⥿��k�Ue�z]ݺ�D#=�Q���8�%������V�U"���'#�J���t/ �Ȇ/����(&0�N�O�v�뛔)R��,-��Q瀷���Sk^���+L$��Cg��Z��?�8��=�G�<C(��*9�6It�����f_'�R�X�
e���fU�s�����F�w�qq�r �?�c�
Cx���!+�T��&D��01?2�����AT��c���B��4,y[�W��d�z�]����5�7��P �����$F���l�h��_o���޹q]��&�u~��p�s\׿Wju���D�	�-�U�$U�v��:�S ��dQ?R���C���?��d�tǼf�k�dx�OG�Z���Ne�P�^���J��.49S��ϐ�}�j{�Ex��K0[�cc�r�a�j7�G<���A��������8�Y_e��o�����������"*����ٶB%�wd�hc���ܙ�0-(�h��Q/��ȯ�a��0B���li�Ib���J,�aX7�)�[�-�]$������l�vxc�����F����D	zH-}u��A�w����'�*0��&Жé�T(�8��_9��.�5�q��N�v+�|˼=�(�;�_�ȉh"��r� �X�tV{G��C�9��u�Azw;�v�b0�����TVT&t%a�uj�x"X�y�X[�����R���~3`�/���,��>�P'���B|�̀��[W�C8�
#np��&�*���t��4�[��&��^���*���=� �z�gpȩ�c�+��Gr��-�_�ZE��M���`1e�Z+S�
� �'Ȥ�X��] X�����N��Ld��?�ި�U����x4?�� G��ac��?vZ�aZ�n�q�n�t��Ch<�f�����e�f�)�+��>*�\Xj���ZΏ{��>����[y`��h��J�¼W\�]M~�ȵ]�б�c3%E&#S����z!E� ���λ�݃��!X�wr�<V�l��Z���d��KN�`%�§z�!�� ���fv7k�����(
R"O��Ȅ2���/$��	�W��+�6&IFE�d-|�B����:Tx��,ދ�J�������B�`
�?^� Ӄ&�
/ {M���)�:D��&�B��K�����&@�H��G-���H��z��d��S�x��oU2�-��%-Ν���݈��䃤7I絕�uq�5�M[�G9C4�E~,k�?OLu�yj�Ksy���렬��������|�}�[
�Ï������Z��U���?�	'�'��Y����^X�x���']2�"\e2y�y�yǘB\�%_%���~^U@���{�8�Рdk8�['��TS=�4�V�+n*�U��勓�#�:Ǌ��K�K��kI�T}���4S���g�;0`�����C	=���]!M��V�]��|X��1ب׈_]��I�2�P�uR�*F���6M�A��+ˬd�D!�f|�B�����;W	B�[��:+4�T��#��1I�I|l����<�,�j�*�G1��<��{��\��se(�f˰�Z�ギ-FV�jro`�ڜ�w$Ԫ��Y3|��4�4`�l�)���2�ŨS[ͯΔ���4.�{	�J���<�>u�gR+�����q�%T���N躥p�^�{}|z�!�*#�����vF� �-Ӽ��g�c~U��(yvj�7���]_��x�b�ռ�h����9���>�e����nGf��|��C�&����:�@$��!��H���Z��y15$UE�L�w+\�;k�I��QttOT�+����G�RRU*�J�e���٩�X)�;��iv�W.��
�"L��)w+�r�$k��r�-�r&����})iI�]�ڒ��h���F��(�c[�۸iW ���4A���B����W9�2�/��c|��W�+y0@l��Dn��~8n�a���3Ocm�^�^;�n��:�� ]{�*{�%ln#�m�x{���(ɧ�4;Rd�ڦy8��f ~�6�[a���T#"�<�S�$Irj�q�IͰw�z���-�wrY}��Ǌ������x�2q���c�i=zQhw�>?�$�����b��_��3_�䍁GP@*�C{D��k�9Cp��H�9� ̺�܃,U���1[�jN��&�|��#zumD3�����Y��&����Q�h�n㔚��[~�!�=��+[&�<$U��v���Y��g'~
�"�!���� 5zLO����"�N�E�Wp���F�-o�ʒ	�u˷^Zn*�mɼ��\�]�����.��V��OCE���Y��V4T�;{H��d��'N�A_�>S6N�����8��.�tM�+"�DS/���k��Y�&���b_����SUGeo�:pe2�;�����A��mǂ_�ͤ	"� f���LzW���k*~�9�4�M9vm��Ux��E-Ю4x�̱e��ϥW�@F�d0pd�hn����ˇD_]$n�r���F��t�R�y��|��&�~�.�e���0�u剴�I��������b�EEB���Z���da�LYkDԝ�����<T�g��ؘ�Ki��o�E����@��VS��kG�h��л�7��q�/��9i��ܤ#�Q��
|C"U����Z�����ld��i�8���0I����fQ;q��%�! ��
��Ya꧃�Ʒ����DK��@ x+�"0��
�x�fɶ���2��Y+�F�ƹ�Ӟ��Kl���	�>Ц�z�$����C: ��b�-Wk��B �>���^߰P�y��6�����4�%��O�$CN�*���]�j�G��I���,���¹��i��"��k�*���O�L���$����N����O
�Z�)X�Ev��m�RTg�W����`�0S/�y�]���h��nGB���'踻%�B��΢�47&��A�ɜ����b���!�>��(��#z�z����p<��GǓ���c?���_��W��Q��j"�Zj1�M2�w){-��z�ʛ鵋����rZ��u�h'��P]Z�ݥ���q ��7"P��	j'Ϟ����n����X���A��y��vV⭁s