��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{hi��7	G�����|��4/���YEs��Q��H�9e���ϒ��(��t�.�?�ѩ<�Փ�<�Evj���T�����B�ݰ7� ػ�3��p�����D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[���۰/Zu�(�l�N
nk�����'��m�n�뛗�mF�觴��F���(�wNE)�U��i�ع�MyS���#7���g�/ AXW�,D8lɗ��+�")�P��L��niIY����x��zt<�^��Domq�ّ0DYH���ｔ�����-*��BJ���Y�A��8��K�E�0;Z� �0������-$�ɀ_�nJ��X�F������;�H�'�mb�և��uW=��#ю�@|�5F/�[�R{��S$���I(2k"�"��$��q��x�z�P�m��4��i�i�e��F�llU����Y!e`e�>��~yL��ͥ|�6��n~x8S�[`gT����"y�3�V�&��k-�'�S���TN�6j���^_z
(�0�Chf��Qx��D*�.R;�V��Co=N�%��!T��߮K�1��ʜE�W �<$�+Lp�N(��V��	�2��8s

�=�[�T����k@���L�0j���Ӓ��}�K�2O�V�W���Q�X��}����K���i��P���aF��=W�%�Z�7���RI���1Ǥ08�'W�P��~�b�(ޣ~���@��TF��^c��Y&=挝fm
�=�1��Vd��;!��p�a1�#QU��s
�ߧ���6k�S���3L����^�<�U։ ɬ�@H� Cq��|:>a��r�� ^>�Y��<\���K�*�����Y��#fV*���'�BL��LE�p�~�o������E�-q�H(�B�����b�V#�@мcvi馗{H���!��P�:��(ߡ�N�_�ѥ��Nh��o����EٴQwc���N��G+̮�W�t�"�/N���w�b�ƺm�%��n�d_�C�f5��2 �!��=�����a��&�����֊fA�]�&~w-���;�a�܎�a�m�x�. c�-� (@�����}��fD^��&|�˗ �F��Tn�N,{�T`�v��7�v7Eb���*S[��u��3'�`|whs��';���R��3F�ZӎU���c�e��@q���x����g�/�:���D�\�Z�a�L�a��K�������o�"��Ŭ$u��e+T�3~20�𐤨-�f�y�l�?_��s|��G;	0!e�]\s�;e� � ����QI�����t�i� ��_�.n��,�}�V_-�!��f��ۚT�='=m�+=FH�UP��X%��Q��oP�%
�f�� ���ַM�Pb�,i��.X�ȣ���BJXLS���H�h+
4�8Eƙ����vy}-� ��=���d��f��R���n)�o0�����^D���$��7zl����w�v�s�9��r����������^<�.�|l��M]���\\}�-&��n��e�I�bY�	���Z����6 }ʝ�#7�,�f�e&LBȟ�����.S���8�p)��~��\7D.�m�,t��t ���7jP�5n�az[��I�K?!�԰�:VcA��h�����3 #�t����w����O���E���H��:�!jf@_��N]�[�va��.NT
��?���f3s�2X�6+��o��z[R��m2�����xG����j��E�i���G��	�\�c(xz;F��b�q�~��y��A9��̢(���E�Z�a|!e�q���j�$4@\�Z��nY[��b����y8�G��]t�NS��0��{��L\[��`�ȓ����R�M���@uVe��4=�Xh�O6�!ȅ<�5i<�����`���d3�;��4̰�gp�PxTG���o�= ޼oy�˱w%[��I�+���n���J1�� Ru�i#5�Afv�-��9�w��q�?֘�>���ƾ�~�M'���a�O�����S)� �<��Ԭ-%�.3z�2������Ɓ�r�����ǸX�@Ƭ��yֿfZ������#O�S�~[�P[XXFy�=/����=Ǉ�I#
^��_�Oӂ��
S ���n0�?C��i�c�K���B^�A�l}N����:�W+��?�+�i�Y�B=�n����Q����{��5<{�� mk��_�,,��Q�ZFa�s�h��g�_�#e +��x��-Z͉1 z������KSPz6r;m�:s�t�7��V���zպï��w��ȶ t��'�~�;�.�e�Ṵ:�&�n�BD�tln�%Ӗ�w���
%<�#ʃ��V_��~���ȝh�t���Fh/�!3��2�2�O���D�_A�3����^�1$p���x]z,>�9�ȯ�J���nh�V������}>a|tcϏ	��.1R4��^�|�s�i�#�Nz�'?�ۨi�)�bO�&���R�Y� �$ԡ�� �Rծ���>����j&��@3�Sƞ[m�ET(��y�c��a�4� �q{�ߜH�C��|�ԍ����7�\Ep���[�A��?���I"����u8>.���6buT2M>]�v����JYW���[�_f�v�=��?#LB����l���n��k�0���40,�b�Z쮩՘���8�0���)ʡky�	M��-�U�b�B��pc�� w�mz Լ(�p�/<���5�s�t���Ҙn�4|�]���(�^��Y�ә����]�f���ڝ���ת��09x
r}��$�T6��߯$_��)��A� �������v�Ɍ��3�7�4)�2o'��s|ɑR��g���� 1�gY���>���%Z��*Z)���/�=�K�Q�B+�	e�����\$�*t��@g���{(Иu�c���L&`g��~$sļRL�J��$I�(��.��ޮsi͓8D�2�?6�j)�)j7����y���[7y�C���$�5[�RD�fT��.w���%�O��N{=R܇y�_�~n9T����M;��� U��U�ī�{Ѩ)GJ�|B9���!�#!'o�������,�}���N/�z$Cx�%Ao���p��E.�/��\��{P���)
���`%�����4��i�b�Fܣ�Ck��f�ƕvp�#�*��w���rVI��B��$oG[?�V���m�Eyx��\���=����x����}�	U�?�(i��z��Kt|������'���B�ڃ�@��֣xkN���e��]E���^�x�ߒ�c����|�q�yƟ~r��L)��Z4��C�l�~wR����u��l���Ҍ�FW�֟�P�"(�LJ�gK�@iL+��	x_��EmZjC)�������/�+���_�/	<N/#e�\m�p�G�&DkK���"f�\|�] P�,�<L[�Β&r8�V�Zp�ʥ`j��<Oe�͑3����r��:����f���ʝP��7/K�86m"J�ɜ3������ns�`A5hn�[��as�q�DH�UWH�����S���?R��d�V�$��^��>I�^>�H8��,�DH+ux0Y��pδ��D>�\T\5�7�Y@��E�?�0�n��h�)���L���R�8ajG	隃	e�x��Z�X�����j�0��mn�U)�-�v����������	�t���{B�}*��#���_��,38�sgp�UB��d)�b���H��Y5�]��=CD0�㩻"�r�C�0���?*��-����Yy�g6�|���)�xC��8�-������g�T;4�L�Z����x�e�wڃ�h��vjt�0a�B�h�>|��"a��&�u���ÂQ�#�z;\�A\b��a󆄧EI�98�;G���uX&�����ɪs�%Yzzj8�^�{}�M64XJ�j0I)6��i1�%r\�y�-��"�n���^��E���ً�!��p���0������ȫj��|vS�>cE "1��_g�������rʄ1�,��rzΒf���@���[�F9��h��E>/�wlb,26����J���%����37z�����1�-H`ة1��H@���|鑴MEU�-��ј\�z@(����w#?}�C�\���"��ƻ�ճl63��������rWx��:�IԤhv�{�7��T�WьT}_o�0`gQE�x��_�IWv�����9����S���ݡ\�k��?7�,ç�=KB�'���{�xO�5�\!ď���\}�* ��ޕ�@/�/N�C�6�jv��&�w���G`J�n1{=jYX�o�����1�?>=:���Xm��+�󻡛N6�f�am�	�������f�W/��Pk��硼�菐�%$p@���"�\���;� �Gw�#qX�(�.�x�|k=�nT:ki�B��.�ʠD� �AeB:��=��Z�I6��'a��6{�;���r3�
`����ǋ�b��ykj4��g=guą2�ka��{��`<��&��zU�*Ŷ9�gv��赼����H.w7b+a}n[K����G����Ǒ�q�m�m��5e�h�9O-��o�]%C�6�5��6WWp��13����C���O���2M�"��,<r��m{�K3��8d�},�ֈ��~��*�ى���ۿ��r��Y+�uA�� ����ϒX�w�M�!JJ�A��E2K0r�L�u�|�c��_� ��On�F��^�[�,z�ή[�W�؋�	���?q@��B��+����r��������,GI�k�������T�� x$�O�Q�+���L��k�6�6Ͽp�H��{�����(yk�m�h1�	�9�W��XB��
���.�v)-��砞-��/�D������a���O����x��^sU	����a�$�"6th��a�- ����^��@��"��b�LmM �	�e>���c]c�>���\[0�a�9٩���m�}��m�DC#��S_ū�I�"�|2�e ��3��9ͦ�����p*���������,X9��W��[3��$l3!��Yg'o}IP���{���H��GK�&��cH�]�X��ͭk���᭝ru'<�Z��cG�S+�g���^��A
����t4A�
<#�r��ԋ:�et�D��e�U�!M^zZ����Ƀ�^\[B��sUSzG��a úZ4B�%ھ�j��-�(ʼ{Ȗ��r���SF�a�,�:/6\^�x�{�(��+�Mk(�5�8f=M�a�(�������"a�ޱ:ŋ����u�J� ��`�5�#��F�-��L�W8�5'Z�S ��p�8/��,ay"x�����R�4�&n0Q~�um�s�ƠM���t�Q�:_렅]���J�����I;�_\�X�zu�>$��"S	�@ �n�3����yq�hX�Z�]R?}�O���נ��OƝK&��X\��]�]K%k��h;�A��R-��}V�)�=v'�ڴ�Sc,>�F��Yװ�-�\e��f6�P~��%D�eZ+W��_Y�Bt~*��pO�_����by��c�5�̀I��J���r��k'ҧ������D9���W03�t��e���G��>7=[![DD���9]}k�b�����zS"I�b;�g�'�~�Vx��|��שFڢ�Ȁ�P��7��j��L��Jz�5�\�S��7\ �F�Z[�d.�F��KhJ�H{xF��[>��IrL�#�{����Ѫ�yX1�x�n;a	�����xƿ�y���W�x����'���h��B���P�"V8D
�-zՅO��/���xQ���B�|Éh"���Tp��s�j�$ב(f*������3��9a��Bb0Sqo�n/t�5Q<��i�����/��QG�d�^@��(��D��|=�4�tu��}Xx���L�����[[\P��E�\ǯ�BְI��V��R�<�A�Rͥ�J �\ā@�b�j��G���TD�
�.�[���_-c�j�þ/�_T#;�"m+M�_����Yb"gCLP�b��i�a��4�Z$�ο�X�|*;1�Y ��{�4*wږU��M�*n�XLQ�3���%qq�-��D� ��_ʏ�C�����&�8���+��� ��|�:x[:�>��Iًs;N)%�k7r�؛�u^ P�������}e�����|l{(�!g�&�{�	���*�[��V�d4�pJ�u�v!ܣ�mLP~]]$�O���,_O�"Ԑ'�ٛ��l5F�O�u��$��E��vN���[�(4?^ _��2N>H�*/��J+e��s!�Hd|6h-	��-=�o��:s��~��"&x�~PLc:�OҟK@�(��=~���&�>�_���4��UeN����:�J����-R�`[.�$ͪZ֣�N5Ex,݅��^�b���k�\h�~{_��nX��-F\����TO����S8����;�?�Ea��0<�~h�T����!Y8�!z���چ��[ �\� �yo��q��>*���G0�ת��qLboE�)"��ZOW婺D�����VN��n2S��T/�W�v,2s��C�~��0�^D�G��lXɉ2@����D_--7��e��+�nP��Naiߡ$w���+��'Ow�J�J�����s��
S���Wtrn�����mksDEy
����"��.��T0pZ�!�!���K*:���G�	��=d��AE�K��� �R��.EM,�v￞Z�I<�w�uz���y���DމP١e��RF���\R�?|U$���7�%&�iS=�XvЀ�:�Q�y��G	9�Zt�Y=#CMn	ʘ�/�4a]O0sg�p�V�2u��z�J����s&=),�]�n�h)9�Ε`�;Q�K�� �%��hU�D�Y��	G�+N�)���M_h֌�d{ӻȅ�Y��-��)ݦ����UܮW+t��)ߟ'\{�-��4W����ܵ��G_*!��99b����U�7�3_Pt�(%�ߕ�6�k��$#�r�0N��J��bˢ���Z��w�$qd3�9v��wi���<�@���|�d�N�����'���l����	�ɕ��X��Q�Un-�}� ���)�rԠ�,��C牓8q����r��TND��h��E�.��J릘C�~8�s��+���|�";6������Њ�e|�q�>tW�:*+d��D�.:^+U�-�Q,��d�g�F&�D<B{�g'$���82!w�2GY�i:�)���Қ'1�ݤ�yy�C�j:��K��6�k*p�uO63ӂ7w�w4��:��;oÜIA]�K��[��1�{�
p�%�LJ\�	㯤ŧֲͅ�
�^|� �l7i����ToxKh���i-���6�n~���3j�	Vd?p�p�շ��tأY܎��20KYh��_h?t]��=#y"���"�wC����j4x��I�@&8POf�4������^���ł�\�LPC��ȼ�����qu�ʙx�LB+{��Ȗ=�Fڭ�#\[@����N~WW��ɏ �v�'�Z�����-Z4tJ�C��l�1K4��K��e\�9�_�>#�k�kg��T�A"�-�6z�qy?V)�-�s�<��U�G���j�~ѻ�$}���x*�[�c
LҖ�3\ �(�B�h���GF�����2ѳb9���")�(>E9"Grd�yNC7����1���E]G���:U�j�ͬ���=�Px����w!3�E�Ƿ�5{4���H��l�U�z����m=U��W,��6�\k}�1,9lq���tb�w�������Ҭ��*%"M��~��hO�D���eE'=�W6%��6�M��/�#��x&�<-ݓr���E#��)$ eo	0p*l*WGi�ܣ�ϯN��L���+�����"1ǐ?�u$5�S�|�u26gaB�ߎ��G��B����U,3��n�+8`Aa6����a���=n,�����8�J�g�X-��-��m��A�G�&��A���w�W[��(�TZR�b<��7��r守 -�EWN�	�@I4F7O��,s�� ��'vv?���:� ���~w�AyDթ�2-V�ԃ�S�9t��*��+A�;����ΎѰ��=_�ͦ7��!�K���h����)�kO�\7K�N7�G7O�	���&b3*�=�0���@�yZ9E�����#xſ�b'�܁y�˿�� �H�r�~	� �4�7�F�
V��c�<�&S���l�\�c �#�O��ɾM.���l M��3:�*VvN֟�������i�#&2=.u��($��3g�+�zQZ\�|T�¼P���"�κ�L�3��LO��;�b��`���
� ���Oʜ�k*�g���(2��5&�seiN0��]�8��`R.���k?G1�gd�"k��'8���P�oP�f����|ǖ������>s��Ȓp��
��&N����-k	[X�(�H��Z´�i�q��~��i���/��v]
���a-fҵ�F4�om�&�v�ߔ%�y��	]:�����bj�
o��K7_�����u�J�*Ğ�ͯ�"��@�Bsl,�
p���^WR�O*U]����f���>�jS #%�]���h�ʓ
ݿX]6-k߻4H��˹-��)T�י�6�L}��\)� K�E�d� �?�;�fg��_�'8����1823`[6�A@D�����u��g��A,�MԵb�7��;��L�3@���ǔ�5�iU�eq�]��]/�����l��t����{?m>��	��D!�\��S5x>���4�+WK��@�UiP��$�޽�e�A�+
��~�9��z�;Xb�ܯ��s���h����c���`���)dx�
�n���W�L8|����k��D��X�8�)�>2V�
a�w����7e�ѥ�d:�׿"�~��?��%�B�����ߑ*ZT�#�O[�O���|9�:8�g������K������(Tpg��u*�����0��Jְ�~���t�L*�ׅ�C}��R�.BZ�n�������y��Ȝ����`�t\d;��EH�fj3��k ���"�5��Md��	&��J�2ϛif�~^d[~ �Wm��:��s;�]b�ڈ����+�k����WV�n�ԫ n?��%��q}�@��z�X��RG�ւ��k�1-e��ڮ�(��@�]N��'/��f��a�.6Wa��*.��`��Ӷd�^i?���ú�M�l�֩]��ch�L�1Ʉ$�	{��R����.|�N��������l���?�=i�T!��O��ыL��:��YRa����|�	N�~.^2(��Of3��L�ʷ�c'�:��I@��n_R�\�^���	��ܾz��n��n+Nrm�� ΐ>�}�E�ք+��:���4D�����򸩃��7�FR��Y�q��7�
�Ո�p�2���,���H�X�Ϳ0��W�m�6c�@������K��� h��� ��L�	�R���W�5�U;s��4捒�#T��Z6�|����/4΄�,��7ޞ����%dT�2�6��5,�,���o�He#�VBS�?Y�=H�I�sE��ڋ~^��,��"�P2�޴0hÿJ+%�`��U$�Xo\�����
���� �\�wsu:��]	���GÍ��&E�`Kx!�gt�L�3�]1f�|\熘����M�2�#��'`����F�ʯ+���~���^�1RL�Z03��,Y+~���4�RU������A�u�����6!0�D�E>�4H&'s��V7�_��0�#.0�8d.�:�=�Bq
�M7`ۑ^���I��,rCa�
��d�j�]������]P��&5���ط~��f]0�K��Kp�<�ۜ����} ñ�c
Wx�D|b�[?$<��D�t縹���s�oYl�JG�������bA\\�'T�CM���e9.>7o��T�ه�"R��d'�\��7n�=���D�7�>$H|�ڸ��F�Lb'pO�o�V	�֡����Z��z"s��Ex]�u�[H�#�kVQU�P�-}3�.�l7#5��-'���y@L:�jn�<Q�'gk��g�$[�⸊��\��x�_2�8�ǳ���Q=a�̿%|�OCl:��iN͖a9��F,�K����
G���v�|B����;-1^uՑ��	��F�0�i;��輌"�n�iQ�� (�DtHG!�,Ѷ�5�o
��֞֫oz7=�����9���Sh!�x��P������t�����-4j�RT�ʄ�����������9��=�W���a6�R�g3��ԏ�����_7�0���[,�n)��kM+[f�UzmH�Q�P�e�0]����Pi��[o\��6����N׳j���,@ʷZ땕��t���*��@�2�M�[�)��,t�����Kx�Y̟���>H�ܘR\��V"d�^�_pm��K����H	@ǌBn%�ê�n����������^�uοSi��
�0�Z����fs�/���]�拒t�޵�R��ɺY4n�7��?�ݲ�4á,ԇ��|BS35�Ȉ"@x�t{�*�d~�_azG��Y7+#��XaQ���)f1���]1(��a"�8��:�HV��EH.�����-URN������Χ4�ג�����br����>���2Y��c ��	]/~�X�hx}Lo��o��^ӏM�kZh�d�GO+&Pu�g�?�*�G���n!������K�G�Tݏ������9�t=�/J1���D�	�ηx��gK�7��1��5�wƯ�{���^�����kVz����#0,�"��f��7�i^,���k ��F0�Y&�(i0�3'7�3���IT30�Apiv���:F'L���TGe�9i\zŏE�>2�m(F�ru��+�t��,�y��F9*m��	"~!֘�Mq:c���g�[$)�R�	���*��(�<�O�N��8�.eZ�-�]M��K��Fi0Ŧ���ͤD�LO�ۦq��\�Bx��RK('�,�I4/�����%k����V����+p�UoWM�dR�&��F!ߏ�<K�[?�٦Ya�B7n�F��Ai����:�^��@�m�N��I���/ܫה�#�j���	+#���.l+q��"A�� �*�KI݌�y��f,a� S����=��1��ުC����;K@�X�m%�h�}4>˹��Ӕ�z��	9�6g<s�ò~�1 ~��y�GY��v*����'�I�k��qd��[���l¶����ۀ~+F�[O��&?����3�b�״���@v�@K��"�'��îh+�����X���"Lo�Ő���B�s�9���6�ky� ����ϐ�3��Q�h�e:��u����|��s%)����2(���ک�>r�z8��W-���ٯI���e*��xs[�HL�l�X+S�A!do&��ѳ甎DF��@vAM�D�K�c����?�~v�ϕ �H�@�������`^�Z��x�cn��Jb�������d�e�WW�����4��\&��aV��A1}~��j�_��"ag���!=Ov� e�A��4S�z�T���;#��P� hE�g�V}Ǚ	�0��7��W�B��Y���vM`d�D���f�Kj�a��*N�b?���5k6�a��M���.�L�ǯ]3���9V�I����y�{ʸU�ڪ,�,��V�*[�eZ��������2y�s]�:�[6=:s}A���
z�B��W�XC�]�����D�0WG�D��05��9� �@܁�D�J�����RA.i[s�(�=?��C�a�~qw!A��T<��d�T�|"Qd�8��5�~��I�Y�n�&V���ňx	D��d�q/�Ӵl�h�R=�t�J-����q�i6rz�/7Ym r���uJ�!��<!�^;W̯=?�����;vH:3���T�R����"�R�fC���+�|*��3�\�+&���}~����FVZ^8{�N)�[#B��lˢ)J����o�d�I���1��X�&|B_�sz�\����eVl$\^��EщQ�w��
e��5�'����9y�6U&s�Ή`v	�֩㪥�{&g��M�jt��N���B�Co���><K��L�<%+�Zz��K��^�Y�l��4�\��Xԙ���P��A���*[��W���g�S8)�
�Z<2��K�/���/?0% �Mdګg��R�o�1Q[��7:����E��`e�Ʈ�]� wg\����W��<fۍ�g��<&��Sr�H�{2i�p�2Ԙ\�.�8`�a�I�YE��6P}޷x�$+g�{鲏����7(��,pO �Z}UbsɟjEj��H�'�v��I@Rr��}1I����]�H�W%}�$����QJX� p?���䈏���K�����O�h8l��]�	�yp�-�U��2x�|� ���]���X��'!W2�x������5��>�O8_��IU�%�.�Jr�I��i�x�%���Oq�-������_�\��XǄv��qoŁ��U��7��fw�jhō=0$-@��U�����q�e�.c��'qL�b��,A���U_O���~g�A��r0w�ג6�����w`|����gm���#��tVI8٫"�բ��}�;x�?�x�#��և�%ط�������W��	ɘ��mb����aJ�W��e��
8y�1���3��5�P�#�L"8�IdP(����_���+c�|��lF �(4	����4vט35�A���qA�E+����n�I��_�;4"�i\ɴ���(�<���Ps�/_��>&B{p!1�/	�#'�ow@���}�W�!+�d
i:R�& ���;`�����n�ڹ��ڿK��4Xk�+ր�?a������S�^Jgp{&��k`�ĳ���#��qQ��:�@�$R��(�|7�ʪ��W��?��@��ॉ�x����}Ɯ�zv<f�<�h�K/�=�%c<�~�b1}���	,2>J���~�䢈/͎^�%V{������	��]���(0D��L�ґzN����%���ǵ=��G�nZg��:lwD��iŊC��W����¦}�Y]���a��r�'�	+dR}=F�[��\-¡-� ^>O��p`2�/v��ڜAk0�(zxǎ� ��㛂jJ�09l6�,2���j�R�3�o�.+�.֐����T� ̮1��ah*�.@��a-��j��C� |Xt)2Ms�Jn����ޗ�!��r�X"~e�c������@�c���d]{�ۏan�0H Us�&�[����c�U�����ҍ��f��dL'�Ø\Mw-Gj�@*�}]0��t����ql��=Zd�GX
A<#g�W� �����Qb�s{aD%6��✚P�Sc��ED�h�܋-bf��|�C��i�ⰕNN	Z����	��A��Y���Zw��h��o:�c�ǠaI �$�?Z���>�0]OGCd �ũ�O��ٌwJ� ��7�q�3�g$
�H�?���]b!H0yL�ML$�=�I�I����� �D#8��q.b���٤��P�uK �L/l�޾n6�bF�ڡrЃ*ub)���z�#@w�alSc�>���PRI�	���䐲�o���q�U'�łݺ:�K��ԯE<vv�O����;��^�����3
M��9�k�L��ڣ�gʖC�Q��p���S�X���5���
��h	j'����ѣ	�[��+=��^�[�{��С��<�k�2D�F�hۖu]����T��[t��EC1D�'7B}� �)pcq`���ʾn����O,��~��G�=��^W��5��Mj,�}��~g��gn��EQ&X���k��G#^`�*��T�]Y�Up�*'��Aд�l1������r@Vy����Ϲ�#D��r�����X&�_��O��ly�x80w�u�<��ЋZ�U�QxT ��ےQ�L;����<	[ΓF{�y��o�qw�By�$�a�%&Xs!����m��礆Eb��	��>T��h���9g��� sΗ\��T3a���٦%O���9r������裷�R�;B�X��`�8<�D�sp�d_$��o�/��ؼ✜�ltQF�5f������S��g�g�9���"�pv뛵�ŢH;��Ghq�l걲���~e"�:��7^�Ļ�V1mH�օyN���P���Q��yj�-�C��m��c7B��;�����;0��Ho����R�����?�c0�y�˗�U�o����� ��\2y���ݹ��#;��Z�G͸���ׄ���7���Γ3�Tu����F��λ�^˼��ޏʃR��V�J�%�S�#S�U��#m-8��?8'wz'�w���<}Fv�֨�c�:@�yΌb%:�1����E$�R��_�%Q�}��� ��` D�,.��Q�f~�`� ���23�����u,�N���1��"���Ws���Se�Ud��EƮH*,Ֆ��֣��G/G֫pu��fD�ruv;2���J?����E�ݘ�B6w ��[5� �P�ax�������=DN~���G�y FN����B��< �v��0I8l�D4��\0s�]���Vm݋N��+��bY������w�Q�1�"Q �qq+�-�'��
��������b� �HaBf��&C�<�|��2��:����� ;o�R�G�#�hg��'7��EN�z����<[�n�^��j7�����Gr1�M�Zȗel�e����Z7lHBy/^U��}Ƌ;���� �l�~��%c�����u/qy��+5���)�@d�ܨ�ߘ(�y�5��g��Mހ����G��_����*,��m��CV�I�f� ^˟%ฃ?H�g�#~b��k$X�ܶ��QP���f��?���wd:�H8�ւlU����.	�԰��SC"y+kƮy��V��<؎π���*���p�e���� ��+z�#c�A��@)|�{�Q��ְA���e�|UD0@��K	�,F�^�E���Xc�^kT&k����e�[��I+P{ә�j������ֽaJ�1�� Կ���zn��S����:M��t̮�a�&9��^w��v�&"/�pE�b�Wޝ@k�<� ���HĀ�}i
k_4ϙݧatβ�����ks�����,�0�"�p�<��%]�R�0V)���a���7� ����GU�}����O�O�'B�N!=�[��{�yd'�%���l�A=z� *A�B>����qHԯ\�S(`�C���n�0��xPj#��<N�I�v��w#fck��@<�;������b,��G�:�r%+� |�4ө��z�3��ʬ�9���4�ͨ'�0U�fkǌ�����/[�!$���U���o�G���$�6x������̂!�<�n���-<��B���v�P%�W�5c�oT��zgIc���un%컞�H)�Ž�
l` 5MV��0�$�J�t�h�� ꐘw�P�Na�*è�eH_�clJj8��)V�_���QVh�I�s:���:A���=���#�܈�訔Oo#=��%�x'�v]U�i��f����5��L� -5�Z$��L��{��8��g���l}�aaag���}��@{q���(c-q5��.z��x~
s��8�!g��z���BZ�N6kD��x�.3�4̥���1�
����X�;�X�Om��iT���3�!!�
��ٿ�_c)��>`�MV;�}�"'��(v�R�v`��}1��&����lb��� �-U����S3��H�8fB�i������k�	�_�P��E.�k�ב�N���%M<�ba���8į���5s} ��&�!6���[h�'=^��A�]�[K�.��0���g�f������<՜Qv#'ZuyROf $8�=�fޕ�k�����N��7��p[$�)E��=�PF��K���^��BOS����ͮ�A<
$I{�hpZ� (�ӈ�^�e���϶L|=P�p�y�"��<��Oi�
��r<�Ozܥ�0�����}�����?.nke�C�c�󵗎F?,Ī���<�������{�/�z�x��#��б�?�Ӥ�rr�����H�l���,I�Pk�TE�8�|f b۵`=�uv�C[����b=���Sůf��,����,�].�1�F��	3cH�ѹ�Lfԫt��/��{�e�ޏo��v4qP�$w�� �zK��P�L��7���X���m�cO�v�g�����t��{�Ւ�����?�0&��M�_ʯ�-�0K+�ԩ�� �6�N��e�k��CY��-fZ�G�p(ۦ�(|Zhχ��=�|*��Y�Jh�>��]�T݁�z�r��K�O���$�C���F�^p��]5�	d���ΓO5��W%���Ɇ7�ri��5� �l��)z�.$�����u��m|}��L��^=��vп�i�02�+���)�[2�3�h�R���7~�I`}��ț��I8��S|�e6d��a��#`N�W���Ry"D��8�j��DX�_�	O���C�!��z�)E3�O�.Q6pA�Ni#����n��U��р}h~�u9r?P�U�p]��wd��/ڳ��i7��z�2��xƉ���G@*�ꘓ��f�Z9`�w5����%�6���\8:���Jǐ3O�ږ�L}���'�/"������`K�x��Nz��,�ˬ�c~<����%đ��|a�j�d�^�A��p7��5Z�kw%8m���x�R8�;��(�55 E��XLK��NC{E}t���`��G���UW�as�d�4JMcY������R4��~�'��[�a�`jׯ&����S���ܿJk���f�s�i�$���&]�����B�(-oԢ���N���y������tA���7�s�J+P&�?�2@�p:�5p��2�H�?D�wM�U�K�y9�#�[�.�}�`LU�0��5pJW~WO���H˖���n�@|�7�*��R������Xة��ޒ�T��J�ݤ余�_Kq �û3'���[`�8�Ֆ���_�3R�ePaS�	�W"ݦ}j��»�5��͕��;z����8a���ɏ٦�5�^7�%�>~[�iCžʄrKWG��4N�!�[�n�Pq!T���~|�j�mRǦn���_ʀk�>��֫���!��9�f�vg��"����P�h߄�yx-��cʙ'e8e���A��	�up���Yt8�f�~S�n��d 3��x;&{����m{��q�$�P.r���tC�'��˟jQ�>���������Zh�:���#CS��6��%V	:��Rk�(En~<��:S��!׍>����
��]1��(-^�%L��d��U� 5�ʸ�J��:D�Fs�3b:q��c��r��<V6k =����-�9�7ww�5Ӝ�&g~��`�p�aU�Q��W�P28����k�d��3Ȇ�������PX@�br��k�YYە�[��C��xR���w�l·}atSV�YUw��/�1���Pc�A�f���C7Q]Y͌E����U�;�뻿�O�a���&HX�
9�0�_�-��g[����8F9��?Φ&��=�I!��mix�i�TDj61P����L{���n�jEF�U
��e�L�Ȭ��cwne|�+�@� �m���5�Ī+�)/$#�"'�N��?�-�F��:B�\$�fۄ��o��Q�e��y�%�}�%$Q�d�rCjxE�0��%���6K��_�QbB�R1b(n�{0q�qu�6�78�Φ��0Kl�$GuO����ge���u�fb��r�����[���K��pb��ߺ
lŬ`t��YQx�X�b�Y]��(���[G�6x>y�	l�B�j{B�A�XU�$�H��aQH�iY��h3Ԥ��B�d#t�{��H�֌�+ӸI�$��+�x-�ϜՅ_ym��X�}���qo�$�~��"��<!nŻ	��;�M���/EB�R�,)V���)�i�/�v8?b�7/�p��C�Ny�i23M����y$6��B������i���tR��%��­����"�Q��j�*2���R��s2.ax�1�n��x�sl�bE$��a����N;v�J�}���ئ$�4Kk�;4v9Q�vj�>�}��X���;�(��j2e�=�l�r��I%�'Ji&w�`�#j߰�K���l�\$!/U�/R�@C���E���ri/��.I��Q�pyOG�.�=���L֡h�
�F����ޞ2�V���GG�/|QW��<��QY}'����tU�p����t���p?mU�3�B��oӸ�)9� ��F�ƀ���~y<�V�,H��_�ĤkפǑ'�����D��V9�#��s�R�O ��O��RSTq�i�4�y�F�N3���)~禈�Nr�G��1˱D��N�pr���,qs&Ï�_CS9z�+cL��`]��]`§�f?���a�}T����0fJ��S"���i��Y�'�i��U��6�?�~��LՇ��Rd���?�bG�X_#�sٜ��" �甡%�}�mM���9y�OW��{��bh����B�4� �$�zӂpi��;�_8?��G�w)��ߧ���T<\� D��t�32��(��� ��_t{������J��� \1�]sCW��B)f�����y�HH�%��X��q@���`�-B���-�j2�8x̛�o2���3e�d�իE�pb�QǼ��)��
_��!;OX�,,��SO��M���2+]	ViP:�R�чH���Z��9y���c�5�$f۹�Q����L;������~�!a�/�1u�������n.���yCz�B����� ���]M��|5V�%'i̍�����c6�0g��|����۰�[6�f��ըy��DJuc��ū��:΄��ҏ�u/x�����ͨ�2ԦdȈ�>�`#�ṗV<-`y��$��~b)���1i����pv�ɸ�������r�h�(S�~^�w�ɈhF���zǜҴ6ߴo���Wm)��9�G��WvV�S�]�2��	"O�: �<1��<u��S��K����������gE#��J����aM|�����G8@�(��	_�{��Ɏ���4�#@��N��)��?Qݻ����N���5{���@0��!1��Yd~��o�Q�1���-��jl��N��+�\�wo�C�*��g�!���8���a���12����Y!��#m�c��ur�}/a���?S@4��W���w{��1}ʒD�*9��?���FX���m�<�듅��"[Wg&��h�3��G2��wGPc�5�t�VN!�K֙�BH��N��(^Y��: ����h\JY\
���Ǭ!���w!B��|0�y�˯ �-oΚ��b�Np� q���L�<��I1;�Ϥ�pS΀9n��菐�7h�C9�7���g��ݴ�O���r���)zɁ��Ɂ���߬ ���^6Qj���w���}�`��a3RY�)\K/��a��W>���^#����&���L�M�Ke�κG{��E�q����#AY+]>�!"�)b4<�|�0"n�����h���\�%07�}cٔf��6.$�����<��+7Ǫ�+�7�i���n<�Cc�鈁�z_�w�����\�T~�o���)_'6�W��t�{!��t�ݍza�7W��a�J��v(���gN�1U5�mit>�:H<�	�s�*jikH�r$�<>��r��u 6�C�;-
"�u$�PrE�f�L�����W���=_�Rbv�����}cN� )�Nw7��91F�o"е�& �3aPy/p�V�?��<��l'gTԓ��@:
�O�_Ft�n{�x"��^t,��V��N,~b����l/��yI���8i�A�O�-�^[��u'����N���۹�s!#�lZ^��K�~�>��Q*���uI㹋��:cAG�Z6�.:��ׂ�B��t�*B�';;2�J P�����_w$Hn� N�D�7$࠿}���tL{�q�޶i�Ĝ��t�J/���N>��ҳ���)B�ѹ�����r�0%WS��蟵^��=����^.2b;8�j��^��0A��g&J�Mo7✒��SvK�K�5���N4)'��]ɦ��ʨ@��+������2���|C�vK��ɴ��cz�B��ET�d�L(pu>_�4߿G�t�=66ʟ�mq�Z����,K�� �����\��/������S01F��C24�� ?��i� �L`�[��N�h�J�l�Eկq0��So
E��fu�w+1�I��u�Еp/<R��i�D�g��]���S��S���feb[�Z=I�Y�e=;7R��"�$]��5ML�.,�u}"�C<E�����n���ajY��:iLҨ(��c�~�k;����>}����ś������#k�{�6�c㪪��2�WW��GcHn�wN���%��m@l�k���&/t��[��6dn�~%2o��U�H͘�+���>����'U�����Hn����۰}NE��Z�pQP8�*{O�b��vq&�~���)"ǧ\��B�\���H����w$J m�z�������+���
Z���u�����ёf�$@�h/x�=g���	
�(�w`��b|.M��?����Zk+��W�l�5��Z@ �F¥��#B�:$���A:I�l�N�ѭ��ز�%Y�Wc
C�=�()�×,�����uo��+��ϼ�8���x�S�[��C�L�^�
'�`�nމ%����� ��'���+�q9�B��,��7#�)k�>�r���LzЄJ]��{�0nv,οi���2��K`RV1��n�,z�;�"=t�}���h�w�su����?��c&�>R�<7(�D�܃�!�"�El�!�pe#&,��;�H���2���6�r�����#���0�á8�F�]�Y��Ut�Ϛ{y��Z	�#�4A�֨x˶�t46��k��̰�T�e˹hh���W�nf:>��^����(�0��E6>vR�N,���ƌ(�ab;ic�9��o���ǝJ^h�t�F=���uf��R_��l1�����Q����$Xu4��H�n��Bzu����=���6,�?]�y�����\��i�~���q��*�f�Sy��]��f@�[8�/�*�}��<�q�.U�ŗ�����J��:�Y��
.4O�$��p�l�nW=�{�;юx�'�6��?H�ae���!��جpO��{�-W�S��D�v5����N'M�O�<;�b0�ӝU��!����QV0�����fYN��r�:�0�G���?��+`(���7vl���|��/Pv�3��|��o�;H_�#0.(u�̉�+����26m���B�Rf��[.�n����(�cD���R#��Y��b5g�8�#��$+�����|#��uWzӪ��
�^�-����B��0�e1@��|�{�܀��^�f%G"�=��q�y��������2���׉p��=Zx|4�`m,�i�.U_Y	:�͔yO�P1�¹�!�:D��?5{�ŌM�JhH<�|!��F
ñv�ӇWO�0���L���quEXu�/�O����44"p��Ȁ�kG��*(JZ����c�)�-�� x8R�m�(#�è���X%���t$c�7  �ͱ�\c�s���^r*�њ�U�r�މ�ɗ��?�o��t��_�����q���-�{=����E��{B�R�e�p�ے\�Lq2�7E�/��tx=ߙ��9t'�8�'퀡�K,k^Vm��X�nu��ߒY��VO5�V��b_�u�+N3KE���"^,�u;u���a;4WB9������In�)零�rSr=R��?�9����Ю�j�`�}�$ռ;�)�O�\��1���h�x�l�ٴDf��Q��j�D2������"�wKf��S�}��g���6E��$T� �Fdǎ�>6l+ ����\�H��.���|'�VM3��|�B���]d����D--B	M8�p1DQ�Ǡ�h`���HU�'G/��	m^U���@(�gk*�:�(���b�z��Kh1�`z���q(A�����=�˄=V��1�e��~�:��N�r휞���y��~����g�_����AU�����(3�s��!���%�k��ΔB2'��5}���J����/�z.�+L���$�J���K�8��9XΘ!�N��x��3'��x�����b"�F�m�w�:�Гq;���0M�ϸs��G��uDi���A>���"�er)Z5�̓�ym��	��B*ﴘUE|Qt�4�O�ݰ��f��6�#�����0/���{����l���bR�{�T~�T����Sk�&���i��@�ACj#�`�
`�������gm��"�P���fU�d,��א�NǼc&�"��~Z�L�r��
߱�⏻��*�IG11��ȍ�0.��r��63���T���r�δ�Y'- ��������l�S8T<T015�8Y5F����)u8���jm0fX�>�p;��4k�>0��&�0�خA"Q7�Ò^��z��:;`����N���""k������R��>�4��2�w/���/�(3�`���d���J���O��ɞ_3H{���I��`;'�:�Y��3]pT��/{�k�#�Q����E���=����҆�\v�
W*z��u@lC0��.����]$�������B���@��g3������I�ު0e%����X�&��R��'�W�%��)��f[LYS�X��F�tn�Ms��9��|��̪���j7{rgucǜ��[�S�6ERG!a��	2M�s�d���
���}������ﳊ�����Z��r���v���͜�ih~�D/�"����<f�zN���70�-X��>-�����(,#�_�����,\�ѳ����}qd�ְ�zӭw+��f`��b�c|v�X�:�c��_�5'�"(=�ӕ�[9^zP�&����Bo�/�����ƫ���Z�C�Ċ��]a>T���y��cZK.BJ�Z�Hxu'^���Y��X�vh$�!�ķ�����i��#�/�8����S�P�	�są�{k�{$�������z@��}U�^qRM.U�Pщ�
\q�!��6�0~0O74�G�6�Wq3V�웁�
�w����aދp����%{��^����ˑ���X0��������v����7O����Gf�z����,��6���R�Ё4���cQĔt.؞f���h�����fT۱�EYr���^�]�%Ƽݑe|��x�8~�4F�.[�^J��.���p�h�j�A6�0,~��q?5��R�h�	 4Yg!�_��(f�@g��h��#8t9Q��Q��x�T�x���a7�i��T��`+�.Wes�<Y�F�U���#� ր��6+�h��
TU�F�B>���&m^�����B��{H5	�<p�iu����4����1>}͜a��z�)�e�֦����6u��Hr�M/k�� ���w���R�Q���:&W��JTp@`��*2��F���g���&���
z�"�Em��ì�GvI⃿��8sת���;�	��0l�M��s�����\ޞO� x����Q>�ę�Ȟ43��^r���Z�'��[x"��Q��'�F�0���?qx�n�YOX���/A��<�~���9K���6t���+��5�j"��9�)�r���T��Z =�y�q�7����q��D~�k�!`+ʅP�m��8,2�+�hL��u~���A�eүE�F�y,��x�e���G.�b{b"��|YDw���\5��'�>X�|�^����"�o7��0.��
�+��r�ݟܸ���*p�Ty�3��.A/sLXԾ���b�c������ĳߛZ��;}.�s��=��̈U(mm�a���� �Awu@����ó�����uMQ�;�q����ws��:$<j�
����?���w��tuD���:@hi�r�߽\�$z1{�F�z;�y�����ϭ��q෨��ɝ�I�/`�2�����6��z�|YJȯR���A|�����
;������GZ�K������,��ㄩ2
H����"����Y��z�~\��v��/oZ�p�:]�"P��5^������K�'�0?�5��e�-=F��>�=�;�L��� ���$��E����.�lz�2�s�RUN�Gܩ� sF��оT1'���"��"T����1�X�ܬ3���f��a��JX�O43e��4�z^ip�;�>�E�YA�3�.e<G��"�O0�
��{�1�<��1�QA��S�S��Դ輛L��
�y�sF�V��;8uS�0 ��= �9]5��	�Bt[�Q�F���IZ���K;P%�t6�]��!C����d�d��̮�rL+yg��2����0�B���r)Nn�!���;�@5��*�N�,�'�
�/S���N�F����I4�Pqv�$�ى-�o�D��0�8�۝�G��H����Ä֧җ���qI���3!��#+�fi[�f�=*��4��_�[��-	�R�J�q�Py�iΜ�'��/���F
��W�#!J��!��e3ւ���:����#^FDN�'r�R��1R:I9�8���C��m-��!X�:�xԮ�s/w�Α��Y3��G�Yȣ�gK��e#�!\��Μsl���'�S��4�U�P]U��2A�( |܊�,�'��c����}��(�"+�%ܶ=�Y`��ќ͓�7	������<vLm���m���W|��JW�O�{g�#	4�����@^�k�I͓<7��}��L�<��&�Ǖ���S]k��\�Tn#���Z����*�^����>��x/ز�K\#�J?��r?E9Vb\@f�����Lü��9�l3��������|�=�K|`?�S0�����#�S��w��;�������~���Q�o�V��4S�a��zm��Q!�w�(�Ƭ��Y�N�FjC �[#�%"ɷe��G��b�w�H��'��]%+��S9����P(�����i��=u1z���\�h�d�`&9/4sK�i#�)X�`�!�z��>��* �6_���ȕ�Kfڻؿ0��幾X~��d��~���Oϖf	�TK��x�)|Wb����h6)�/��| !�����E��6ƴ��k���R�����ؤ�z�R��5��z�P갘 3�m�8�����8/�0[HsN��%��r���ד���X�h���~�}��?W/���X�N���~c��� �?��v��b���Sט�U�)+�͔:�������6��F��p�	��|
�AQ���LU5��÷�#sG�2���z��W%��� Ԯ�s��3tR���0p��vì:�z���͑�'XvV?IxA�I%��Y�a_������h���9|J�U��IR����dXچh2F������˅R�%��X��`�sf����:^2M�N5�ƚ�����;�;,�`��Y�&�b�A9�j�8���EY�/AZN2��V��	���40q�]w�����e�؞
�0�����~".*�����-rKjrUKk��ӑ��Xd���!9�Թ�~�;s���CԧO�	�����_�����e�j��!4��f�}
tQ��]�7F(�c���1Uk��j�!�n�H"�6�(��N�ħ���ԯ͋���.`���w�Ճ|�)-�N<X��K,��6w��o���<��jR���@c����̈J�`'�(W���2��)Jk2{&0T�'v�6% \�>�����J���|�Z�䷥����gȁ"خjO�#�n���k/,JZgz��O�t��}z����S"��eT��ۉjŌ����}�R��@	��҈�j�Q��¡V�5]#K�
�l,��� 7R��U��m�p�R���"�\�<���o=Xui5_��?�����Q���N;���ɹf�B��
�q�p���R.d���1��}	��Y�F��bKe�c>.^E�
��٥����!b�~5t4�j+YlsJM�j��8_�����m�u��'YM �<"�-��'�rRI���1��gl^p�V)�a$�#��$��J�*��]�K�xFD����6����u
�(�q��\J�p�� ]��Q[A�
炴� ���q"3���pzs���G�q(�$����V�o^�ٸ�#S�D�*�Zxs S�m�޽�L3�eX��b;���"R@n%<X3��ׇ��V��F3�?mc�g��5���!k0�D��#�CQ��gSq�q��_p0�E��Nָ��D���t�~�_,�^�.��16���w���D���Nݽ���T���E��������_+#�5�A���c�LF��x��?�nL���Qc�&_�v�yFF���:Dۅ&�IH��s��嵏d:�B,�6"�{^�F7e�ࣛ�e���Ӳ���|���!BKH����e�vָ�&m�����þp�5ۙgp&�j��̯������Ǖ���[���e:�Ǒ�{���ϸ���ց'1$����������(S�z��o�EEGVƾ�!`�K�a��}Fj⾡�Ȼ��ꢝ&�x韐��د�I*���=��۸��o�@2�fI0��V�����e�a����)|�Zr�b��^��\i�^�]ߔ���3�.�l�D7F,�5�7ɚ���6u�o�FŤ6�g����E
Ĉs�H�ɊZ�uK�r}�:�6�4Q0�8�qq��eJ͚�ld�y��0��E��8 �eM��G4�Y��, ����;��ʿ��F:��g�P��,���7�j� ���*ίd~䙕�o�9����K�e�+�iK�>9����b���N_1kZ�oO!���ٹ$3�7UB�NA��><$m}�����3���Nw)6I�ZM���K3�}���xYL%���D�1'�߮�w�������ḟ�r�e��p(h����_W$2R1���%�Vn���U�R�Ww�v3)�����2��BO�7� ���--��?�x��tSP�u$.b'�|mrl!���W0��C�-�} Iq���;��N�{OiO��Ln�NӉH�y�2�� ��߉w0E��W�+��w��=�����4��
u���1C�bZn3��B��y��O��Ry�6ʶ�G]�Q�*J��� ^qĮ�=�D��C3[^��r�h��5|�h/ѓ�\�/�w�s<�_�	�.J'� ��/���:p*�p.x�r����,���E��;20��Tj����sFB`�1S�o���\w�i���;Yh�,��a��G�6�\�b��#af�h��a��<�Dj��/е�0Ψ}R�g���{��*�|7���JD�����������/�w}��d!k���DTz@;MP�����(} �v�P`u�/+Gv��<-O�=kf���Ē H�t�;�V�4��D��B���|�-��6���9�;��)Ϭ�B��Q�O5Z���q"��#��}R�"���/᮱��nY '�~�¦ H���c*�}+Ȧ㲆���B���z��I���m����|d���)��8��V	���[�C�}uU��N	v�i	p�.�c�%N��JXY4�0���
��^��-�+b���]�3����#�fT��vb .PW�(���<!��E�#avQ���ߌ^����� `���p��ӌw*��Ŕm7h�@��_1�=�X��"���d�ޗٗ#��(�a�����~{t��p<:;�W��bZgp��p�LT�گ�-�����fǞa�Ã��_��Q/���`'�Z���;vZv������6���	ן;�z�Sb���3|P��y���!oOD�D�]�.�p������m��kF�F�!؁��H:sA�x��{ګU@n��y�QB�/j�4����;\��ʘ����v ���"�p�K5����y�.)��g���F�Q;Yy�TGb ��P�3��η�M�~oh�2�]��{:�y�4��V�^m�ː[� M�T��ʾ�2��%t�3�Ju�a�� #ͯ��Fp�Z���{��K3�u�z|\����#\^�:���_�"��������>��tI�����G�b�_Dd��F���9�#7�Q)=�D?çF�-

2# %�:����O\�/_���S����>N��'}�E��gf$҆����"2�i��(�J���,���c���5���Kc�W�j�d�J�%0i���}�~��#���;;Ī;���D[ڴp�((�(���M�x[��ײ��|Jcf+{޹-C�m�[��G��v'�9��ᑔy��sĮ��%��uy$��Ay�[;�,B�8���;�Z��PTl`�q��p������!�z��(=5#��|�����-�!�&�O�Ӧ��9����i@��Y���
�08鮻d�+�O�yP�&Ꝏ��2>A��l:=��.3I��5{S%�ƁM #��%ml��:�kuJ�p{@&k�I��yξ��- ���MċD��_5�u�� U�_�_�e�� &E�8>H/�N�d�U�$�`��0H�H�'�������מxk����}I�o��1�tps�6�+%���9<lb����I؞9�D��p��+e�=�7�[GX��o>�<�?�RNz�gLYy��'~U.������/zx'�s3��n*�^j�\-��9c;���y�D�ba��G��}r�u��ƅ!eG�B��4�m�����i�ئ�ʤ��^C�Y�7��7��ר~��8��ߖaY�gn���\i���g��=�7�@M�싑���^L�_�_�-�='[9�
�k����V��O8*�&Iv���)����]_���B-x�Yx�
���y7�'S� ad��P�ɻ�������_�_���3w�K�$�j�w�|JSg��?%�0Q#���q�#�~�|:�/�RC�.ס1Ʉpl�aZ9/�g3T6��H |颅�qԿ�rt]�*��hW�[��I�.EwH�L����uy�`�%�3�ϐ�SMu�wޕ ��m��W��$�]�U�������K��W�x>A۰;��X(*t���bTkJu7��f�d�|�M�?#�z�ݘQ���1�@7�ƛ?�QdH7�O�P�!X��e��*��7f��9�|�wh���sF}p����3�"�/��nX�vGHOS���HF����0���������9G��}��G�g/�A
«y��_��|*W/�0{�^*������.�'��z�oM΀D����GEʾ����mR�N�kl������i�L��#�V�C�N��`>!����M����u�6������P��0�{^83♀�vB��5lY�����i��4�mr��ϓ����Q�"$�|�n��c�J4��e��^� 6��iO�[�)�$�*��g���E���um���dmӽd�.��eݹ<�=�ӆ ��/�gtP����6�����*�p��	��=���L�S�Y��g�6!�U�7�m��S�`jǬ��F�d߱���Ș����k�4���k����w��>�8N,��}��z)%z�����J�*}�6�(����p�񫙩��i��R@Ά�.	��Q��k��&RVܣ�X�M7�����a2�4��1��۟�5-�_e�u`��ŚF_���V�W��+e=�g�|22s�1�l���2�7�_DɎ�L;�����P��w�ӆ���ĔrT��j��OHV�=o8��F�ܧA������L��֙����3�Vۤ�	C�`�t6B�r�������A�L���B_��祳��BB���)��Q^�f0�d6}�-�L����b����D��Ä<Uoix6� hE��Ma��wa���Y��͐�vX�s�~���ȡ2�K�����{���RvMw�RBg(����M��|XW7�U������2.U�h7f�I$���C˶�ZO�lJ\�^�d1L��n����K,0��ק!TB����\��4�?������x��.K�������@([���T|
2��;�0�s4��q3L�����x�XIl���g�0�ȋ?���� m�5ܹ�ң��i<��8�]���VP7u|\���9��DG;d��8��\���I��ѭ,���po���h=SC���ۨ�@�a�������YS�p
��l4d��q
�i�<j��VJ2#�I�E�������9�up0R�x��?�:Y���@��aI�A�	N�q��1$����\�q�y^�́D�3��J�ߤ�!`�L�Z,ѽVB��|Paw�a�	Ԅ�\U/I`�w.��/���L� �)��a_=��{5ɗ{��7-}�<7T��Y���!o:�� ��e�wit	��|�Xo]��&�ZÝ���L(k?��W���	.�ջ��&t���V�@7^B'�xj��ܨ �vޱ��m d�$���apN@V90g��
�k��e���w.��i�qDF��L�V*V~P%�K9��5�\zz�J}�ڿ����s�b��~1��_]u(��;���1�V}�D���N�Q�"����&j%� *v*���
x�ǘ����8�_�ĹR��c