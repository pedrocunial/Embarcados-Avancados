��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cЦhUd0*$;,#���iI�2��~�y�ܩ�v�iN�	u��h��d�#�,y�=��̌(m��B�	X�"�[m����#�邂�1��F��i��\v%h~��$�R��b��b��Uzs+�>�<�i�������cQ���Lt�b����h��zy��]A���gF�ŭF��~�B��V���d�}W�[�Z '�B��@��P�o�C�>����z���=:v"ǜL�ܬ#b1x�q��6�±�5桖�A��
"Kk�:�A�[�u�;���e�ԥ��W����Kt�2xB��~T�C�@y�.
_���%�~�d�U�c�#���E���	���E��{��'�L!�+���c~* *��ڀy5���N�GX��?�x\0x6<�<r��˴�8���0`�Y��r.��*m���X$U�ae�:��
&E�nO�I#VŅ��i-"���������w�D�0:���2�����^��4;�2ǂ�ۆ�M&?�'�%�@�<uS��r(�cԹi�O�cgX����a������f�>R�C�l|�tD�v�"i~=�0� m�%||dfGn�e�\06�M@�Ѡ�V������ꈝK��gv����/C@�=�"���m��)�cM����DR���\��n���l�j���A���#���Ks?�B�Roӆ���^�M�8D�e��w�y�0c���S48����q�3n��c��.���4X�:	5T�q��΀>}: "�?(e��ВQM��=Pǅ����8��=>m�d
�N��<�����Bфj�ͯ
`|�[>���T
-D�=	�9����!4Mw��������e�n�ٟ�9)��ֹ��l
�bD��F"qQ��H���kK=��� ��!~8z	
 /�x[�8� ��t�(�0&[C�ȅߞA�:�a�133�0�I4��K�̭�z�Sx��#� P�ca�`��:BLI���ى<�Y���c�]�������YK��Z*����\�o���C
�����^T�rE�^%r�>���̩�)Ȭk��ˑj�*Z}�ns�!Q�O7'{n�k��=~`��ad2$�q !�\�(���l�cMpz�ars楬Rs���W��f� �=�
��/g.� :�-��r>/�Xm�Z˥v��8�A�$���֠=�#w�vK�����MD�~GW�^Ň��o�b��S=���6�a�\�O�t8j�ת��R5/0J�3�$L�;Yٻ`���4|~<���Fx� H��2���|�M�6)�7�R*qVs��f����L�n��޺��^];dB�ch��b�gMf&1�X�W���|�;�ܤ��ʀ]�a){�nԭ)m4q�RA)����kRT�3�|(�"n��ùŻ�hu׻�o���m\!���/g��͉�9�'W��v�?~�=h��ɮ!�as�cZ>�@����5Ͼ ~��J}8�Re�N~4�Z��;T�����9!���r��ۻ���A@�X����LhY�]�F�N�&'Q�ǭU����âD�ߤ[E��c�q��C�R)f�%'�wyG�t�A������	��z#��&��11�#)��P�b`n~^�po�!W���/�qV��@�̰��po����3�_?�8����a�Yg �I6��w9��e"��6�p�!� �i��қ�k��1�p��>�aA;���۰@)ĕuOS.��.��X���	X�	/�E�轑p��.���0���Iۿu5^��<@�41��lŶ��,%t�KR���8�I`��$0�r�{" �>^��]�'��o�����v�>�3e�+��9�����DHr�d��i�x�"n�dK���(m��,��e�)��|���D6��H��{����G1����F��Z0M$ r!��ǒ���(�����K^��a/ �O��̃O>"}H�xo_&B��g�,Ս��Тr�/�(�d�b��;���5!!6�uwM�P��j����S������[2x����2��M�-���v�!�@[Xv-�:fIC`N`xɝ|��,����rGl)*��.�lh�0��~|e�Qڗ��Q@����X!��[z�������+��"~�:r�+���^mâm���
���1޲��^
|�.�?�<�]�1�A��7{����H�<&�ʪ���_B�5�vI�K2̂��5LU���r@�g DxSx[G��J�i�&[P9�5N[�Lk/͝<e �&����_����=3�z��m��{=�u�H��$�ޚ	���@o�4+xH���� ש��h�br����=����\릊��X��������vGZ5N�<�n�R���L��-���zC�!2B��$9m��5N_ԇ^.�V�{g�S��6��%`�4)�oiO󉢉M��#��-]]}��|繱ƹKNM'EԋQ�����	�Dފ��,��?���m�3�X���Ϸ��t!�I�F"w%�O(�Q*��c�p
��:�RXF���s:(,�&�o��		I~���&ȍ<�㩙����-��F�Uj�����r]8�AlRӯ������g�@����_�)��\%��6E��K���m��P��W����}�9�BM�����j<B��zQ�h��.I�g|�Ėy" ^�w�D�r���&^����Kb<xD�5�U X�	"EB.b�.�V5�z؈]�R ;+f^����
��<�PpS���<S# ���Ƌ��|ٸ6Y�m!7���ю�!��>�h�ʹ����t@����SH/�B{Uvר�!�׭v�QltZZ��>K'f�����6go9�,if��qW$��x��e���[�������pg��B��L��a�����Tz�v:F�8T }�C�C*9�>�ϧ�q��c~�|����Uu���g���ˑ��3�L5����-���_�,G��@�GsIJ��'��Vz�%���^g�"��Q���;�q��DzL�-/x:��y����h�=�q4�l�O��'Xs爨����B�j�B����
���X��7螊�I��!>�N�,��>�\�y���NA9�b�e����j���MFjg�"?�42��B�#/I�C�+�򴺵���W�_z������W||h��w%��L^�uW��}z��gk��*��R;���qs��&D|��F-�(����Si$:Q	�ڥTmg����TbA����x՜�w�?i58�ok�J8{�̇I��2��[ xwQ@!U.�	�Q�����9e�ϖD��a�4U�)���»s��x�1>ֆ���4܅BSn��6��P�o�\��v
49�,�(�~����JE'�aOϢ� ~==�7SY?Z�c�� U�a��:u'�����Y��0��&Bi�qjƳ�o���b==����{��kK�edu���F���?�K��1P���XӋ�Sȡ�]k��y�7���"u}���Q�Y���j���5����}[��s*�����Bи�"��w�7<w�]5��c����P=���Ck}[��2��&�t�h�{���};���]�B�(� ��Q�/��	��MVM]���<9Md8�D9U���/)����8F��C0�"ԕd�eV�x7b�
�ߌ�Q ��ab��� ����Y���+�E;�R��P��d��~���U��Bt�� ����7"�C����8WDD�2|��ك�m�*s��ni@��T��.��4���a��Ǭx�+�7ȽI��W�A�b�7��כB��p�.��#�k��|\�a>}�s
	`�d9v�{e^�va�jM��/v��\G���mP4��K��e��c�+�V����M��_W/%]�]�H��m�u�MF�趝�>=��:�_�a'�����/�u�f�T/�O������&>%��
2�ӏʒ��
� ˬm}P��Y��w%�0��`c��S�n02���'l��`��)��w�d,�pk.:�oa�d)�	0���_������xs�Cҭ^NѾ�Lk�d��r�|���w��fU����X���,ҲN>�}f.}�\��xL9�NF�	-3 �?�5�6>�s�����;ޑ��}�z����[5el��P�V��u�{Յ��!_�k�m�-'���	�r���Zh¸�)ظ�����#�:��J��W������a+r�ws�}>���uۼٶ�}�Yn`�ă�a�w�r���Z�.5��E�D3l�q�A�y���Ш�ZLOp�u��4�NE;�`{`��DԖ��Y��¢�w��Z��N���l-�]a�8G�
��,T�
���P���ϫk�ɕ~w��e�3;�6�&C�\��8�!��Y(��;=pHT,�A��w�!�p�oq�{�BQK�Z2��l��!�~ڿ�^�ޏ�yvy�]���YM"�|&C�.�թ��O�����&�}Yn�E��3��n�ӆ�GUo���dx���z����y��5z�g�J�B�E�*4'O`��VŹ�;4�	�}�D-i��#i���jx��u�J������ Q=;P+^��ofp�IW(˭=(:R@��˪&r��/ۄX��b���D��P�Jhh�3��t"���r�I�S�h��ԟ�`����r� ��P}�}@�����.͛P��+	����PϵT;����b�)�\��Q�g�M�?��?�Ż�m�o�-]q3��k��
�}�jF�ۣ-	IG�n&�Oh5Z�5�!ݒ�k�����{�1�t��?���*kQ�3����,c⾖�d0���M2o��(�SO֦ʟ���D�]�G�[�q�;����ײK���t?h�(�9@Cs�������!ۼ+�x�6^y\n[��B;Od�T�o�����2\d�� ?�,�7�e@�Ӭ #����+� hH�ϴ�voڋ�Ǽ�����Q\r�-��;�	����`�ooK��Yj|ʂ�{�����!�����8�ՍŜ,�1��6K�q�����ɫ0�Ŗ��y��n ;�4��5�I�9�҈%�o��}�0�Q��J�[���z����l��K䍡��R���#e��9/AS��K���!��5岒�歂�ڣ�_�*�Xl����t4�/�4��+K��5��z�;#	c��n�S� �� UyYl��?/7-�[��a�[pѧ�<98���R��F��}��6�2T�֟n��?3ӡD��������
{Q�)Q
5	K��j�yդ95���g�iصn_�%W�"7AR$���j-�8���́�)F��h�^K����%iw�0~1k8�m-�t
�+����7��2Q@��+�U�gr:gެ�k�oR~>�������`������@�b)# ! �����	���x+������Ԓ2:p�+i"���O�j�g}��Q���3���j���'��3����{�P�/��v��4�+.�(�D����^'�j�W��pυ(��n����?#�������o%��Y�PX�2Kf ����kR�8��2|��u.t��g�2�*K����0D�(�^�F�i��P_�v۶k�;r/P9j�"�� �XK5~�$�U�Ϫc��9��H	ш��z�CW6�"z;}�'�ӫF�F�TM�2�RQ��6 �����D*�1�M"R�$	�i0{�P�&x��ADI���Rtۭ�b�&� ] ���N�XmD"�ԩ��<'Ψ�Ъ��18��Y<��J�t1��%��<����Zo�O�/{�_:�����|	ӁM'�9'���$��y���C� �$3|lEd1�Dvy2Ɇ�'݃�P8��7��u_��~��A3C+ܒ���>�c[��]�I+�[��rq���4�S�<<\`K8��*��1�Pgt�u곒(��r�ZF���36����G�n�K��6`��µ�9h_#t_��$
�An�c���_�g��^޶�D��_�g�6����h�M��n��w!a~=�����/��!^\}���k���}�-W�JF�.�nv#4b����v������F(��B�����YX:P�~�#����|�o� ��=�<xeu1U�bz�Y�k�c�q�Rp�6	��k^�A��tH�:�Fg6-t �0`�:wUn4�?� �tc��YDd�Z��n�Y&�Xt�E�q�W
����2{�&u�#β�j���_�2��<������[ҩµW_i(��M*О��V��\plc1���c6��a�[i�w���$�^0C�%��z�n"�B������wW�B�OjY� ���ܬ'r�"��Ϯ�_	���׺�x_��b掆'� R���1e����|�'���	��u����)� ����sztK��D%�Pp� �2B;Hv �0LA�����-Ƕ�cX���x顅�[@D��@�6��\�G�jp������/,�w�6s�;��H5H�7BB7����[�P@�����f����}|�GB%d��6(��*��Z�ڏZ����P�rp2��O��7Sַ�B��������kqzx�B�rǫg���54��C�Oe<�Y�鯗���9Sr�X\h/�ʖ	V7�k��;����I��T�Sv)�]~���%�
��fq9��l>���Ywq6�WdK{�q\A�B"�
m�O��%�����Z�>D0����8���j��P��q�_C��:�>x�0Ldz(D�R7�Wn\�3�Υ��%n��s���L տ�U����@��8����솲�<�Oi��By�\�%���J�a:��+���d��ɫP�-T�6І"��є��D<k�%{��;N�0���I+�<���]*�׾=&a���(D�>�M�IF"~�\��4�<�v����눮�l�
Cб;�hB=I��y�������j^%f��3A�����6��v���?l�^��	��^�RA��|M0ɏ����y��sU�{`�=Ċ�ϱ,�[�6x9�7���F�ZN��NQ՟��y��Z����ݾ�7o���U�^���/޾�>C��ݖ�el�" ��5Ѳ��:W�8��/��aG xχc�>~{K���5/��G*��L�ĩ&(6X�vơJ /}' G�Eۈ���C>{����Ϊ���{�N:���KR���qλ��f����Jg��ds�ڎ��(�c��lܵ|1� �����@;��8�$*��1v�լ�)�.*���(�h�%f�!O{���$H�1����[���6�ʖz!���<��c���q�*u�������X�W��ĳuv�%��U̦�r��z1�Maf��5*�!^B��8�%��O�g��}3��)9��Q)?Qׄ��A�ػ���#�3�n�4���<�Yd�+�� ��lĺ}&Q�E�xc����Q�o_�6�����jgA�F�謱�09�%�!��� =-�3�81-0@|��k8T]۫�M�EƓ��Ŕ�(�lr�2�W@x�r�܅�n����&2�w�yE.,Uƺp,��&灝�~lyÄZ���ػI@Y?gt�\^0_�S�����h �@������cx(�S��� �fY\	j�x���d+�FD�����%� �ak�z���h�"��p���4w�����g��v$�pG�]��g��k�)Y�D�1��D����<T��!D,4yU�{Eܯ.�0������Y>vϐ�����K��m�,�D�7���O��Χb#�'�'ϾSH���q��(�?�"�Ek��D��ȕ=��ˏ�Q��Pw����[�N-L����ASEв� ��d[��=N�l�@z����TL����?:�\��P�d���I��AƼ��l��ڊTI��y8�$�Պ�cӀ&5Tf��{sՃ�P�"|J/H-"R�=����R��:�/��z��;k�qȯ�
���m$�d(��̏����/�>��M�հҦ�M/���;���['�	��_����ՊBJ�]0p�����������`QO�)���f�����މ~L�d?�Q�-`�I~If��F�f*&����3��Mi7���y�6������S��;�Ht�UI��3e3d��
3m��l }c�d���I�*v�,�_�=���ӆw�ת�3n��Y��IG:��aSvS��?�{�vw� M{ʫ�<�K�J=����gHQ	,5�+�����}��(�7f=��[�'�4�m�a�V��No.�u+"_�;�S3	�x?�N�q/s��S����� �f��G���(l����r�hHW� 쿯�O
����Tƛ|�o�a�Y��tn��Q������P��3���l>D%�bp��,����r�#������e���pe@�y�=��������ː�|���-�����P�(ɀs0�(��#^A��#]�0�!t����5�P����(V�"{��e������t7X�բj�p�Z�L��;p�U�zη��_hdI^lE�S�����$,*_�I�[��R�۳4Н�����^J���"�j�F�x	B з����F��	��hץ7@:�w����q���7z	��:�`q6�J&^�U^�S-��#%��\!��4��強[��&j�n_{�I_9�=�����0*Me)����f3�ݼ<W����gN.�aݕ.:�ޒ���p/p�sW��Ӗl�U�|H��
�#�ယܨ+Q}��s(��JDǳ�ImQ��R�}����/�$���`��]�^�l@���uuohV/�z	s2����"�:�5:�ݜSF����hx��#F~�z�����*�����^��0��;�bO}��}�����{) �)qbvj���d�mm8S��3p���� M]�R����ͯ.D{�/gYku�~olڰ��E�k�8���GCȃ�6R�Z� QLF�L��������Adt���DQ�N0q�#c7��xs Ԇ�l����E ��#�]*KgMOjt��ǔ�)u�� v����Sz�nO�G4�=��02
}�������|+�$��M>�6o�1��}����0�p� �Ա�ˮHn�/���I�#�퟈���V�}[̯��4wy�!��D�JY�hXs�0����]ZsG+�D?�1s��-��a�A�	�qo�ǆ,c_���n] zc�`��R9i�z�O{��-�&��\ ;p�AX��w70]�O��FTp��y���2Mx8�hd3���9�Dq�(4��3~�B��8���4�jϾ����\³T�.8I�-@/�N�H���O�-��t�.\L���d�e)���O�Ĉ<�Uӓ�b"H:��ǒ�-n��;�% ���m?��0��$����5h�?��b♓���To\d����{nu�O�5�潪�W�ud���tG� ��AY�W��7x4C�B�����'栋ob~�C~�l�\��1�#ơ��:��v ���4�l�3�'B�'��y;�O^.��M�=�5��Ì�}�F����>��,M�@wo��`�oZ��I�N�[