��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[���O��T�Bܛ�^�Ό��5i�y�9�U�K��?}��G|��q�v5�@J)���>qFe���5�x�Ӌ�.s=��#7���m�˕1�օ.��4L�9ˑ1g�ǐ�\!8=|.������iQ�z�P��>)�e\�a�C/®^�j�Y�u���8
�5Jw�L7�mC�("��b��wqX,b7��ǁN�j$"��e�)�Hþh|0F�2�_ʏ�:%
��g�R�@� R�~FIM��Y�gz;�� 4�Y�;� ��l�R͒�3  i���<�K���u�Ky�L�<���;�/�f����8OX#�	7Ǥ��@�)��>�1��9@}=ȟlPoc�*ȩ81��$�SY�9��pGy0A�D�[��2gQ�m��~��-�Y��$�k�����ǆ�����M����\aX��._L�D����O��h�D�E�:u,�f������1U���[����O��OS��С��Bd��nX	�7X���Й$ww��ε,�0�O)��¥��W��Aw)4�\���E��h���Vu.��p���aC�Rv��g=cZ�9����0��������;7��w���w�j`Sҗpl��ɣ4�������o�k�/��|Bh��F+��4� 7yq�R�OA>Z�f�'~���\Ziwh'#2Mn��qP<��@��5���1,��c^��ssԃ�:e�7YUt��h��J��^�!���*�Ā�B!�Q�(�}�ϕ���[�6�#�>�>M"���_|�f�Ds������Y^�.�B�t�F�`��Cθ�����E?m�Щٸ�iE���D@-�(l��C�Q�j��S�X*=�`���I��sg�]n",XoGå��ݝ��~�(��O��_g_�0J�+���5Ce�I�D�B ��2ɕ/*�/~j��rE��
E2�s���N��l�ҽ��n4u����:Jb�j��9�Tᇵ~ `�)�Q�>�d�ε�5�o��V��y���]/���pӀ1c@��UʒW���psSl�l�z*B��.��
=�A4�	Hp���m|)]�T�J��I��%s��>���=�~�>�zU�t> �W���/�
�q�*��"Q�a8_��71���t�P)� �X�[nʬ����}%!�ڷZ�O"��30��ty�]�Ħ��S�`�k��'�tu�"6�LƦ��ί�w�5N�b�clj��\s�9L)��'��������Y�o"�4,8�>�C}��"�d�cڥ`s�˷j��0�wˡ��7�����QB���[P����:Z��:H��"�a��8���J*��}��'�Ap(;��K�k���v���|�i��3āG4g�Nɨ7S��=�I��黜$���Z:Z,%F�̟�{
Go[��r�F2��"qI��,�p��8��"�B����+��|�%D�
'�Fr�����n��uk1����N!���\�����sb"�Kl|�{�}ь)-���<��:�'��&Ě"�rlq�39��8W�jى���?8�h7Lwķd�f�����kHJ�bόQ��;�z�ĸ����k����wc�Ȟ[��e���0�@I<8�����N���1K$��řG�Tx"��%;:\�T�3�U��f���BkN�����)��8�Q�OA͉4�ҴQlmtѽ#��� 3��b�-����%fō�߾���cʈ�����r��d���Ɂ��U�q#h�`G�pLL�э�c=)jP�(�.��_��=kF��^�q�U+��{ �W��g�ޖ��&GQv�/�{�f����X��~������i���J�ٱ4c:��!U�	���VʗdyU��+�������nT}]�c�d�o�f�W� �_���o���F�TI�w묽9,L�4?6 ����^c	u.l</��&۸b&�M��@!$@������w	h8�,A6wHL�<��;J�qz9��d>�uR�Z�-K�?�ÅL~Iu���!���ʴ-��1�:�Q��N�^��+�Z����C���Aeo� 0���cA 2��T5B��Ţ��Қ�OBV��o�$�N��?Qfmʿ�D?��k�ŀ۬;�x;K��|���(!��r��u�:6=��BK�=�9��{�ފ[�O0!�n��}�7�yؗ�ܮ�W�������̂�����l_�����Ȇ�2YmϠ�DL)_�D�QK�(+<#�=Obѵ��kn�V\�hȅ��=;�n%-����d�i��7�G�\���>֪��dh��g߈�½�z^N�|��a`!B�č{��;�4��k%������{���_�}��ŉ��N~1��e~,&���XC�'6!j���ݔ�,�#��nS�Pɦ${((�:�\"}�����1T�_�?1����*r�u�麮�����
D�,��'��h�e�d��Z./����=6���6�q$��"x�`B��/$�n��vg�X�95�./����q3'~.��)���¯��S�������%]��Be��ҫ+�3�x�:"�.
VՊ��2O�'X�t���� ��;��J��5�T�τ� ��&׳�)2=
��[�ȇ���d�"�i�IP��Q�4�Q˴O��5�zoy^���P��T���)\�._��_s"=��O��tQ�S��ݢ�#��&�w���f�����+o}�P��"��[�������u�������xX�nM0�\mB��z���a;[��~v\�m��
Aء~JC{�3���D>��,�����4Y��N�LAk����*�M����a>9�U�+�M]nqtE�!k��@�D��`.|۴�&��3[Q|�<ų�Qo�A��sG�ob�2�ĤV�[�h���>��B�n�j�P�iJ擺�#{ѱ�������d�Wڒ|���	MM�e��ۄ���`ۓ;��I���]`�x2:a2KVSrHJ���W��}��
9�r��u#kC8�t��k���+���^��������.��,�'w�<��!T��P)w���#>�`���Nx�Jnuߤq�V�+��c��ؙ�̲:�ʎ�6˘���R�h#�;�h����r=UjX`0f�����msB[s�m��� �A����d�0H�P��j�)���f�2++�������y���|,X�4�;�6j�c�H%'�3��&:�(X2C�X��$�s��>M�5�J��e-_3�K{}�A���qDI���,�<��Si�	�)<��Qo�c&�\/��;��P���˸�)�pJ��h��(�ui��$�	�=�ov�М��VtJ��~_5>��U6��v�Z�{��N}���Ɋ�}Or�a�����7U	+�R���̟��h� K
��"�:!(%T��)".��V�9w���_�Ë�kGE���|d�j][!�G�k����tPK�9�V�j�$�b�ې�ƶɴ�Z��Z*o�|��s>X����9/?tB��Yv�I�h��L�d4�lY��	�|��oֲ�qzO�6g~KS,���H��uI�?t�okk/!��E	D6\`XEf81M��9��0��;S}�t�RZ��ɭQ
�5.�&�v|ə���K��_"O��;�H����8��j҆�0�q�M�ғ��(z�~U����NT��̢����1
�1���7a��	�'��3�˝���<�8|[��I@۫9>D�gY��^id��+i��k]o\�D�2]�#�_8w�ؠؙ����c���> ���a�xaQ}���wj�?_�{%`M�y��#�VA�Q!�K�����d��b	#3�l�{��5�����۶!�}�X~+y?f�E5"�q��E�a
�T-&�6����Kp��H?cI�5k�{��;��ͬ\"ѻ<eW�>6��?,N%�j��8~��H�
Y�dPZ�sV��˄��ހ��� >��"�S�4�a
JuJ�����X�e
�����[�#��0��\rJ*mT���h�[���y&�t$Z���'�0�^AOy�i�� C�33�;�	QO!(����ΒCb��/EjO����(�0�CT���%�<8����Q�מ�A�M~&^3h��%3
{|����/gpd�qP:���*�1�:.b��2����f,��+M���6ɍS�Qj'��qd�BF<[�M�ˬ�»��ڤ�dR�~ �����y>�yMK��L�؜�3ӿ��u�(A���}�VPUŷ;W���2�o��M����aE����F��@_�bF94)��<7(�~];��z�_�a�Ӭ~@��j%[A�n�`&Q�����M�K�x�M�	��&`�/͖��˪�R�@�.w\��
�`NZUo����	�:N�Z+T {v�^"���$/tN����K����5��I�l�`��"3ײ�wB0
ym������8��Z�0�6��r�����x��s��Q�N��y�����u�*I���~���j�ϸ�uH��`+��`���T�Q��aܙ&����Sr#�=�XT���&�K�����6ZF�\b��qo�;_�C|�B&[�J`JS�����l�6�p��@�&<�:�ׅfn�
�l`�u,�v�p�q/tq<������/�@������`�������	)���r�H0�h�8Hh�#�z磵BUs�N�]o��]�����I�t���^�%��s4Vr�?���!�d�x��y{ь6TX;�b�$^�PJ�ze�`^[�A3�*s?\��(�(��P���e���滠��{���%z��}�X�zv�N�5��c[��e�k�d����E�(ã�ǘ��Ԝ���u���	�58��X�4��>1���4#K���þ��X�d�k���[#�BMٳ����"BQ¼��9p�Z�y,�0�g�>*����)88^"=ْ1�m�]���>gL.�{�Y�ne��U��~�� �y�jP5�U�"}mQ���/��+I ��LǇ��"���
�Z�1�Y��{�'<���b�������8F�����~AH}ǩ���m+�c6�W{�.���6΋�y�;�x��J+��Κx:j�|�S\0BMG%�����R����Q����N��q�u4b��U�8C^���58O�Hjo��˦P��գ���f��a��M䣿��:��t�f��0��	m&��u%iKVb��=���g��5����AQh�����(/����H�}�u��ѽaɁ_��+&��TIb�vM�p�6��έ�3;���P�P��(�PX9�H���G2�G�b"Nh��v�=q,�����zw�%�!MD'f���l�J5>ͩj�%\�@�֡�AE1�=:@�(��q"�-vNp[��"_��ϑSw�k���^��E �TF�OPF.8��%z�'d(ty����(���p���"{�k����G�rw�H�E|��E���L�/��RXL����"_�� ���@�{D�[]<YZf)x�<�0��d;�MH%w $O���;��^3�9���ߞ8��,o���)A"��6dO����O">�ځ�ɇ~K��aJ:���56�E3��naG��2L����f�� `d���$ ������J���$�J��$��6�*BfB���%Խ����x��χ^�t��-^$+H�\�K���1_� .�iѬ��jv���?��J�>M����'���� QDەma�#���\���
.���X��J���!v�U<�@�} >�!��>��m<��Է�ڥ���K6�#PP���8|S�*<�G<�Y(�P��!���[�d8���V�F9F�s�4��W_���E�� 4�E�`��e��/0�ļ��v�Oky;���_��N!4n����z0��[ �(�rǱ�H�YHF�e��ׁ��Ɏ��4��k�+'��̹���'�v$v!G�\�q���q�Y�T/⦌Z�����ڶ���-�te������D�9�ɷ=���@���|��|���=/�ec�
�R͜#��� �h�c|g�nu�����i��{���,T��ƎN,&M�\�:�������4\T�M�R��O(-޹s���P*�o^m��z"�C�!ua��k�g�R|uQ��f!�������CQ��d�^���5���*���|�p�� z;��HnG�`ֱ�\F���p�/�QU� ��w�Qn4���'DP���*Q�W�w�e���rO�%�3�	Dʗ[q^1�1򙝞ō���<���P�{X�q�v(<T���&:���/gQ$��F��Q�ܻ ��mX���I�F���3X .���H��?�X�������6Ow��P����_/��F<RTjR�,d��}6;�#؈���b��{4 �|���EAl�O�X�v[͔���'��P� �4�
����C��N�=Um�~)�R�����^'���$��� �Ԝ{ �����Gf��h��Y��YCb�7tjxe�W�'LX=fD���̔CJ����� ���'����cHd�#Q�	�	�l���T�jJڄ7EE��tz���TZ����;���1��I�<�M�2.!�X3�������u!ag���l�$&;A��d��8��M�y�����<�wi�T��S��)�EL�"���т1������B��#��g����`�1�S����PˑΜ��p��ú�'\�
鵷Q�bL�gL3j?D�[�h��r�c����V�\��W����	ћ��<f̍D�wI��d������[��L��`�;��9,��I��V�7�UK%�X��\B7��h&��؏X�S��g��Fpjo����
�������х<���ޘ�DJ��k8�ͺ�4|"n��N�=���}��/M]Ӵ��g �I���>d�$��"[���
�yye t��F�pN�K6�B��A�Fq�3�\W'��.QZ9
��ء	QsD��V�-S��*�5 >X!c{�-g�/�w#{�1,��e��IЇ�3*L�?��[������NA�X�I�~�-p�+���M]�-�1I��-gPN�����³
�Xb�k�	s��?tFܛ �8�`�d;"��-�U���)���`���w:�|����5�i�/R����ސg�_q}��5}��6*���l��l�@M5*������xg�����9���UICҗ��	��"T�bG5����,%�kܨa�h3
���x���r�$�k��v����� j�Tf��Zy1�&�3܆߯���[�6��;�h%�X�@ 8x�U�����Ҥ�t�v��C�8����L���W�u~��\�l/+,��l�ѳB�T�v��T��jr�t�����P*w��;�ce���_�����.L� .r��KOuG{¤�|�P�-���,U�'Z�a1�K�&6��T5���]\�V���l��ӥ��<�/�?���$S�����;`�T�������B�d�X�/�������