��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cЌE���M5o�(��[�Z���YLt�Η����uN�p��K/�p�����Nv���"�ﾴӼ:���{4$]Z�a���.��I_�@���y��@����=���#���P��!Y]O%��sJ�I�T���n�'�&��ϺG(�)3xpu^�7fӓ8��ѢEw����*��!-f��9��D����$���i,5�֗6�_�"h�����⽆��`����X_q��EP�X���H�ͼ��Mݠ�7N^:0:s�c�\��rsb<����| ��D�ȣF�8&�M�^W�v�x�x-�İA]͞��PB#)b������t�'|�~��fp��Y����;�<^�=�� ���
�TfƐ��@;d�D��H�a���:��������<�O6&4�ʀǭ�H�[G� ��^ {q�>��������g�԰D�t�l�pd��8^6��ct7_�<��������80
�����f`�]��bp��L�ma��� �]�C,�oٷD�Z�nQ���;1^�����J�A�	,�3���d}��7Q}�/��1H���s%d�Pe��hs�;�Ծ=:��=m�|���#"� �J�]�k��3��5>%��a9�������MN*�p�s��}��F3�d�J_`�Vit84 �sW�b�1�׺߸>���o���T�Y�
3�����wm@��ՊW��=�
��m�0�h�P~D��I�Z?xɟ����M�37�'���ꜣ)GU��T�+�V�$�c��r�P�ifKC�-�"~q�O�gz$ԟH��c���|���"/��hʦ��?o4܀�)��$R]t(-9������:Wq����qo�<z�-���b��c�cx�V�{$?v�����Q=��Ϣ�p`�A��@�wi���;��guL�{�N�^D؃�'x�.|��-�A�{���L#_��� :\@�bO���i�ߴ��ڵH�Q����#҂���{���?���&˾� �&&H�W�=#Q�Y	!+1��T���a%�,g%D���F�ϽJ�x��Zk�]d����t~+:�|&6��uX�BPd��ㄓ%s�+I	I�z��x�|U_�+��#�>��Dwe��5GM����Y�4�x�,xW3�8�v2�J�*,x4����M'DLN6ڱ�S>-��q�ì���wX��~1�S�o"^���.�������C�D���K��w0�DD��V��P�[Հ� h�ݪHɁ��6%i2O*��$g+�~��`��3f��#�%�D�#���8�-#7|�TI\O��8oW␇Q�8��������"Oc¶H��������-�Rs�?m˭�PԷE��'=l�w�����x�!��
g !�O+,����������C�����w$�_��=�����G�n�_ �5�%��_�����>�z��M����m~��S9�(�_(F��V�K�DQ��s�	��nm�)��ܯ%{1�dVm+�����G.�_�~9"��Bb�ɰR=."V.�u7�./��ɽ���_}�0ϔ��(�>F��"����Ax�K���gl׸ӓ��'���G��
���n��.jF\�
�X��#8ᬦ��|�Jn�0�ȖғmM K̽�v���"��i�y_�6-�)}�Md�f2s���A9���
�Q�R�>�S����9Mj�X;������<6�����hMKk��Ij@?R��c�%��B���7H_��ᄚ�S�%bU��J�����	9�C�!����tvW�u�l槚g�;��俺��o%��nXޒď�ۡ��Q�?�/D�X����f�+�9�Ls�*=N'a�}�Ü�B�^]$�a��` #1��Q����xf2��;6M5�ٮ����0����L�x2�;�ɉ�\2��<��'�X��K�:��˽����h�&�&H��t�@����O��/�D��4��b�Q��d?��a�����R��9�ݾ���u�����Lk��m���Lӎr������)�A��IR���@t��h��m[�O�o�GfLE?Y�"�Ŭ�R^��*�����"�Q�":u$8@�F{MC~+8Tc_�3�r�CJ�ϪFI����_���\�̙s��J��_��/�`����\S�c�'�~�b�x���%y2��|9�9R��j2�Q��'S|B7 ~� ���`гi��0����vj�.g���ߎ��+������~ �GS1�%��A��T��;�;�?�� [�_�v1�/����Ps����_�F�C�w�� 1uAl���	hs�YyS�&�Ɖ��гܥ��*�X�~ح,���.P�V~R����ʐP?d,�gٕ����hV��N��]��{ ��4y�b�T}�߁ƲLSW���= E@n& �	�'v���uܧmR��Z�	���U�[9z��0;�\�o�.l�j�w'	���cxN����1���I�4[�/���Jf�#��g#Q�r�����Z���t���y���O�٧���9�ک��G6??Z�P�ԱG��D3����D���ѭ<�4�9��/F��pK0��BC8l�\4�H7�t��=�B��֥}M�RJ,Ե�E?g�z�ĞDF��LK�fޯ�1��7���W��XF2��'�4ڎ�cJ^����~}o�9��e��G
�JM��ŵ	��1�۠�7����=q4+j�Cy���[3G5G�G׏N
&!���,������W�+S���^)�m:qk��*+"kA\��tUn�ͷＺ�2<�pӳ�m����[�v/C��{����=��0p9��|b�ye�ף�?� �����M���EN�b��>�7lY�X��2���������f;6��2�Mg&㷝��'kƯhz}�I��-�3�3�g���~\�6\��A����������Q,�� �1-����h���1�^�}k��@1W���R�S����Jߢj�%o̸tbf�K�u+Z����9���B,�M���S�C�����k�3G�;�N� u����vs��״�K��w��m���C�������x���a�ȣ���<��������`�d�F�8]�ȊZvcѭ�7��ɤl�_bp`���Bvϫ�Iv��1/M��tZrF���o:c'�\�4Aw����ץg��i:�yՖ�����un:�v$���U9�T�����?�#q��{�cޟ�yPެh܆P��>{"Fm�lv�uF�B˩R�c ���+Fg��u96��:[\b:9@6�V�|ߍ����|�VS��K��R���㏪� ;e�=�Z�"5W�ic�Hy���=:ܹk`^{��W��K�h��o.|�p�8Ne��F���B*|��'me������y�
ReYp�1�/�KK�%K `�90v���mliIs�Nȡ���fl^KNM��g��bd����?��\�F9� 
�Vq�8[���D��(���wg"��J�T�ߏ��z�j���pD��J�'�Bk��6����s(V��5�2�'���fѼ�,@�B�u{�ٹ�e�kּ!�04�"3U��F�/���^Q�J~�|p���w�]�W��Kh@�f^_y)��t9|�,��,�[��&�C=U�&��j|X�!��~���aQg���տV�p�l��z�����G �lbZ��=2�	W��?$+$�����7M��� ��}l�;�H ��ʛAa�&畡�D�$s(Ş�Y�^B�7Ǒ#*f1a.��j3�g(��U��E�?jܤ9F������{�	Q<�m$o���M�#��qF��.[��%k�г��T�I���"A�O��#��k)��E�>���6�3fP\f��j!�פ&X����D�D��mإ"5�K�p&��_�z���H��>?�BRi�S��]7,L�?�ލl��I�uV�Y�"�j'!����ƕ�qA�B�$/X�J��-�$�Yۑ�s��#;��4�O�g�@��m(��k�I��k4X^6ϯ.¨���W�7��g/A��]]U7�S��Z�]����]�	�m�8�2�il������kA��<1�~
�}1j `�iqY	%�_���r����T����K��v�ܛ���S���!G����}[�/�S�Sv������K��_�|���ݥ�Qd���tZ�/��'�Br���G��K˫�i ֒sWX�h�)_���Y�o2 ͉'/��-��-d���A��uv�F�ˈzR�=�)_�1]�*���D] ����5���k<����&#��`?\ݴ�A���+�9��p
|��d%6ӯJW7 /r)��>wp�
˭�W��'-
�@�K)P���p�������ڼ��ݘ:�[���.i�L�`t���6<�=$KԞЄi���S�A�7̀9=������2==��ˡn���c"P�{G���V`�Qީ��z0�����!�2Pz�MKv����=1�rU���W�����D퀶�=��x������%�^��	,�'\���r�H�fc�P|��e�[�q����d�W�N��,���\��6�Ԧz�Z'���-]�h����rB�B+X�Їx���'8�����(��O�������4|��u�^7�I�:������dvi&��F���Pv����I(\1��ʃ�=�W�x}���#A�I�d����>�4�����f�N�R9��?b�W�CDѭ��z"	,���s�8fFg�#�#z^S�s�>.Z���/����G���E7�����S����c�?�'���%,�u�˕Y3q[�����^x�����W4��N���?�CfI*��=�>�4�s԰�Z�`�E��G����X�EWӦ�y� ��w7K�讓g�-R��bi[�i�/�kM�U�1��G@�qDڧ��[7�Ʋѵ<�Ș�P_�SH�T��`~^8��rYV���s�W@2�+F�f�:y�	ʭM��D��8p���\־�OS�X��͛�$OИ��l��ǝw�{���$6EcM$hTs����Cq�[��)Ɂ�ۥ�u�K�
^uK����\���[&<��ܟ^؁�tu(A?�Q}��0c�;�j�`�ǼP�nQc��Dp�I"\@�������T!7����XxѴ_w(}���?kC"�>]����;d̯\u�d�l�����-U�#�"Θ4��L�ӆ�Kȟ���<ȱ��������4kn�i��V�u�f����ҏ��75U�	�4u�'���1�p�";��ג,t�F� 1�Q+'�%��9��ę� )�7zefQb~Kg7Z�	�o�t"(=���Ο�� ;�|h=&l�S� A*��C5��\DS����&��ӍSVOEՅn/^xsG�i��ʖPv�P������%Z��̃�V�g.�EN��,U�3�.��Sm��$`�7avj*��e��Z� �������ZD���i#x�\��bnL0�B������a�_g�o�ic)�:Q��Y,�����Ƀ���{����bF� Yh�ߖs{���y�dSf��'���%��C��
-��z-0��}��V��_��� 9��%�r;���|	(��?Ϗ l����b7��)��1\�S�O)j�C��&#����Ҭ�(�'�:�}FkGh�-վi5,��;�!���U����ڴѲ��&jI6V]rK��'g�(�� q$���T6�Z��{}��>^���1�)a����@س�'��&�?�F���{��&m_��<k�u|-VN��q���5Z��3[�ˠ�g_9Dڳ��ަ���*$��K��ԋ��e	���� ��4K�+���y�C��"�|����u��-�����DR��6q�sԃ�l��f'�����t�: ����.+q������L"�����2�r��9��dc�Mg'˝+lESG"/_"1xh�CVb�]��pͯ��-��hϷ���ﵦO\�K��[�zT�G/�B��>��}G܍In�J�Ԫ[�r��s5%&y�-Ł�@/�u*�6��Z�x��P���}3�*۫C%ݷS�=��iy�g��ؑ��z�yq�iS�8�W^�R���1� �?�S���ȼoD�j��g�:�ڤ�u6��ߴ�^�x�o�H]2C�E�WN���QL�V��8rBI��	��9q�#���8R>v9��O�{��z܍ü3p�5�C5���B0t�����<�#h��A�].ޫ���@&�	*���W�(XWu�$�<u4�O�߃RO�^8�����wI��͸�.�I�_���A�:#!�4F�/�2��_5��s_Mj�
����۔��Тr��� ˽��U�܏�4�k\��Fl�k�*؟a�x�`�߅��J_�$U��j#E��.J'�s3h��"�w�X�p̘d�
7�XTh��{��%7ΛP��,���
tm{��_����9kl���%8��L�иl�J����An3�A�����~�ksÖ�(֞�[��V���\$�k�i�+��y	�P�*���-O��S�@ib9^�EC�L�Ґr���O�xn���I;���{�1	M"���q��<ӏ����*� 2q�����X����hգ�DB����Kfd�x�0o
�Ȅ��H
�c�,��̧�*�hsp� (�L����ț<w�U�O�1%��E�ٵ��Ir�#�m�����Ş؏G���Ąk�U��h~�B��}��8����+;��]ƼDm¤�,\�Ԧw������UhE��A���s.��[�9`�n3�)p
�n3�	��	[`��SْW����BM�o�^��7�3!�s��2�z'D���O�W� .*��x��j�Z�foY>8?^l����J2���B�'���]�Y��Z�;��uH.돇5�ҫF��4<6�wI�)v�)qK3X��v��6#�k����Z'x�HX�5�
�v�%�yh61,q��4�<��ݱ!��>F��)�f�l��K�,Ս7PJN� ��V�x�>�c�yH�5�DY�����sA��:�_�2m) ��=��W!���0�a�_mq � s��T��-�%���#����K���z
��D�Cr*�C�o���%����{GL������I����=Rd"�H�^wQ�1g~'�=���,�ؕsH��1�E��K�X��Ĝ.jH�C�WC����VjZN�� �kߵгhgW��¶�b�*ǳ܈���Л)��
%�F+~�L��Q��V�$ڻ����a���Hr�S�;�v�;�U��Z#��_w"��ˀR��J#�
�����U�W�!��j9��f̰<�M5V���`���s߱]��M���"���{O7���$�\;�R���~��]�m�⻑�L�P����$�v�F�4�ď��b8�	�F��)g�{Btap����^��1@/��ؙ��_������Гo�H.҃T�xtr+xX��z_1�%��yx��~�E�@T���z���%����=�ڢSwgY�s����w�u6�B>>̝$/BM�R�S:T�>����:C���U©�KH<��ω2Ms4W�r�˟&M1�e*�	��d�G�ǅ��2 ����9*]'M��X.�rQrr��a'�G~Ü	��B��4��c�~NB�^��`"�(�L��WͻX��z<�f��˫�z�����.�*�����L_A�W�04]�uǊ���G�V��N�� d�ݑb�NG(��m/�!�dmت��[�����y3��20�<�w��p%�l)�K'ق�>��D�1�ω�[AM��Ӄ06����3r�i�D���bQ-��m�k����4�l.�Ρ_����~1u��.4����Ӓ����ӅHp���\���AG��x�i���X�Qo�p0�{�;Y���6Aᬃ�n>r�|�m^p�
������woWl<���m����6�Nߩ��ʦ.m��n_�#"MýJp����'���1(�A���n۽n��.$�uֽ�&��
�΂U tt��v�Cț�J�UKK�I�կ�����>�L���;��.�Z:q��R@O���L[4�����L�:��j1+r2��v������f�8����OD�����7���}�����:U�-����}g����a�!�;F �(]�O�~nF�d`|�9�7�����V�;F6]=ȉ����8���T��7�b���b<(�n2r��ljn�!(��ا� ̿'
I1�(V���a�>C�Δ��o� �� ڨ�i�/�01��0�A���&�c:��]�3���1(O��ղ� ����8�V,���ܲo�o��Pb����(���Վ��DhӆB�Ր=uCؽrl{W�4E�#�dm�@�o����x�F^���y��U�����	[C��E�q2
��m�"�Փ�"#�g{"���Y��'�>A���~~i�V"12����!x!z�K������H/M����X�&�Ĩ1(����y���X�p��)Im��iN�~}0��^��L��{��B�V��B��3�}3"�D�⓶��I^}|��Հ~�{������a�W�^Mȝ���Sw1�Q��#�dh��1�@�"�^U9C���y=��+�>�s�f�GӒ Ô���s�?�@D������h#����H)$D��K����2������&A��1&���n閛.9�T�r�hț�gJ�#0k���^+`������}�%�����w�:���H�z��G=&Pj��a����7��_���vr�;��Fi�z��٠��̰_��U����%�v{� 1H[�?j�����51�v��\M=�	x�i:a\��� V��8��fgQ�7�����*C-s�f2qQҴA׽���l�¯`o�pY����ę���ǎq���������� ��/p�3�Xd$ӊ��U(0p����h���N(; D�5: 凸��H��͐Į3�e���i?�L�6���أ�S�>��`yk�䫩!"*05��?k��������8x<�&�%�m$��$�󦷴�h2wRTzv�pl���	�i~���4��tIA2��R؃D,��\1��FT����'�`2��������  �c�[��@zC��ѳ�zϮx\�gI��"���k�SW�OlT(�7g�%�	/�=�j}��C�0=�c���ˣ����YQ��(���"��	���]{+JT�}����k�a:�婖zt�R��DS�/���k U�jo�50~��|v�*J�V3�m�1�Q�L�*^���F"S���8O�D�s����Ӯ��z�c*�Sut0��#��e�H�݂��^��q�Թ`��e6Ř�6ΰ�"a;l~���N�pѭ:2� [�(��^�c�mx%,a�%�7����6�!˃I�4{��$��L[�d�Iy����O}�>p5l�
6�bأ���{��//��<o*���q:��Re��K��>�=(�N�4�*��e]pv���e��'>���,�A$��o-x��!;~�\L�r��-�8�j�:�:;ƺ������{�RȃAj��d����GZ���^�j�H*)��4D��0�g�Wν���SN�jza����|}n.�Z�\�U������ɑ���=\w�"*�����1z���!�5�R��#k��k+�G����/��Q?��b�-��\�G�����nm�O�r�ɰh�z�>��'P�3]��tרAM��IM�cε�NMJ�cx����{�w��ZF�(�0`�Tjv�u�K��K��8ڕ_��@7s�暣�DHm�"�Z �;,%h��H����'خI���&�q�|[BR��	�2p����[��۠�Gs�:jt~��g��B�:ډ�mk��tj�Z�~����[�
����6|:��3e��%�z?����Qeam�m���P��z�r�h4�_ 5{eD�7.�]�`@UW��H������~��/~im[�/�ZNS�몀>I
�ZL�T�5��u�9�U{�)~9A��6��\�BN���a{�N�Tb)�¹
���7Q�twو�����T�8��n�<ԓ����#냜�	D��[d����^��) �ѵ��<���?I+��F�>y�3IJ��L�׭����
wJ�4�Q�$rW�	ֆ�^<�z�ٹ�����}����vʄK��*�^[�5�O�I[���V�.�t?�x,��z��R�"���WD��{c�9�5�*�@I�!1�z�\�9rBs���1}�[�~;=o�4GY�T��י�݇>��1��RM�I�K�\�U�0�����
�!��h4�U��vVLnn�@a�2�*�w�{�ݺ�4M�����]*����F��k��IV�D�ҽ�З-�^���F�;�3�Hc��Q!s�G�J>ܷ�`;d<�?���)mH��/�	(W7���X"��p yM,*�Yt�8�x���N��}5ye٧R��1H@4�9d����
O�'/;j~y	*Ə?�)�����R�n�2)���)��g��bt~�ޙb?���#�V8��y�A�=�%}#��'�8��@�KH@���ߔDC�7�j�w滘|���R1�j��*o��z���v1OB�X�
�?N�=wh����e�c�Q�q�C����m��04�z����M@j~�g���T7D:�w}���~:#�w�����6���?�~���ǀ��O8�lG]���Rv6j���fY�:����[\d���KLi�¿#DoG@���a�I��7=��/7��fn���ºԵ������o���@�r��&�(�%��p�
X��(qr�=m����t��'�lJ�+��H?_��|��`��Cg��v��h�0�*�k�t�!�b��_[�����e4���k(X��J��ыY8I�����.���J��.���\A F���DH�4�"��A
~��r����2Y��K�v�{W�y�w� ��R�EdR�ˬ�ŏj�2!��%x��^.�����&�1d��D�ɫ�=��γ��S�=Kެ�-8��n(79]".����q��!m�������:�T�֓-j-oۦ��~��'d���@yX�	�	��2En��Wnnc��\�9��L.-�@TC��u���Յ�Orx >~���HNW��ӕ�$��hI	 E�4�2�N8�^���J�6��G��~"�`]�f���@.ٛ���\8G��"t�*!*9�Y+϶��2��v�i�N+�7�d���k�t�1���pڮ��z��Pk�{�|e�t��9���r`s�|���I��pֻ�<�D����߀��@dv��8)�W��㯡� Ñ5"�#u�.*ݽ���7kf��ZGNݼP���#6��#M�h8=���1y܁A��`�+3H��V��5�C|���zr�jƭE����n_�/�+��
-^��6[�Ѽ�N!r�M�%|���d���
Q�.�)� �m�2�H���3�x-�F��
Wm����ٲ�{!Cb��+�j��Ro��=K��0�.g8��|Y�8�YZ�a���ILYZ����N�(:���V����'I�����k���'�ç�3�(v��#��;���D�^1!	���� 3ɨA��8ys�]�~��^U��
d����}q��$Y���������r[��^�@v���YQ[Aʻ����ł% �s�+��0G�,�!:�V6`z���Lie@���瞁d�j õ���#~����w<FxH�*,��(3&��*[s���N�w4�辛{G��\aiy�)���1����r��=�>�4��1��M6	ȃ8WJNjcZa0�t�E��&*{���_��3[0���u~_|�xW	��;Ƿ��vkW�)�Bp�
=��afs퇽7�s�f��=B )��� ,�O�h�x��/c<�KY�uj`�9b�**�pL�fd�g�ø���u���9�e2h��H%g�T�U��_ꯘ1��=m)-�Q$0O\@�u��:T�#
%D�p:$ѰԚ��5�I�T��v[�5�`�z�Zb."@�p�)k�!���0���1F���"h���E-�S{�F5N�Ű�<	�
��Eף`�����Q!�=܈�H�@��VN&�/���l��
`�t��u�/v8�� N���;T�FQ�z=�`��ݙ��o�YB9�bC�������5�ku�A;�ԛ:ax����d�1�"��E�N��,:q������D�X�n�VFQ��sVWu>в�Q��\¸Ҫ�Ԟ��pn�LJ� ]��#�$|��I��`�i��$�k^�E�6t��@y37sVUM7ݰo�o�" (���!AU��`� �^>nt3U���3��">�����>3��9Pğ&�\��͢f�=� Y}$c1���Bhz44��M�Н�4���W"	p�wfȔ7�~��|_a��[Lb�QG��y����Z&�v�]G��Nb��@�`I�Z`b7o��;���k���n?~!>ŉ�[��k�`{�:�}1�P�ezR,S�}-��_�v���b�I�m�����q��=����#6A١�j�拥���p�0�0�l�k���w��[�8����ֳ��!���W%�:����z��B�h.2�Ƌ�l�8�V�:�BpNكY�s
�YZ^t^.`�+L�I��+(B��Vf��v�8p���yC�ϙ�WU��+d����Є�	�U�r%���r�v��
Io�/���xY������\_]�Y��}~��8�Q�EG��蜵���F��R5�����g��u�x�����L��e���Ƈ�ī��5�b��Ai�N����-��yW��\��:Z�3�x�D:�b6��5`O�I�FįVC�+ү��"�E�}q�E倁�i=��(��J��47�[&~�-J���]���oe�}����g��������8jo�= �Ĉ�5�z��JZR'��i�d��N�3"�N�����O���i�{4�B]�P3��X1�_�UL}�a�&�U�U-#H�H&�#�%V�0��t� Mu�{io���jS	~&˦���F]��_X0X�7�Z3�x?B' ˝�02�)4v]׃���0�y�!�"s�\�����
uel)���3�4����z?0Q�N����đ�MUr�.�x�S*m� g#��qv�A���'=4���d9�q�'��@�x볝�D�!�|�s�	�����	ԛ,7���0W�7��]P
_1���	 ��E��#s����FV��P��&����:w�V�����	Q5�+XJ���X�&�4��M��Ћ^*e�Ͽ�A��+Ӧrހ�6tZ�~�=R�:�dG麢�wQ�E��v� J�)bؓR�U�?���S�y�/p�"�q�2*��p{C1b�BfJMY�'�r��_h(�|O#hïT:�9�����AΣi�|k|Do�hɤi\�Y� ��t�_V��.���T([B���^Ka˨��N�]�;��t�Mo��SYx��}}����X)v�A��ٯ��l��w6K-kk�3re]�!�L^tD��\��̸��\����G���qT`k���K���U[�_\��ŨWK�E��eт��������d����fPnja7�o�O��&iBw��q?��=_�߱ ���Q��V"��u�.�4O�V��=R��q��G�:W�S5��T�TӅ	g�lr���Z���Z�/NO��t|�3^��@��ѧ�>�M��v���7Ea�7�M��vB ���X�"uJi}Pi����x�s�c��tV�:��Z|!��Q8�̕���:�|�%��Gfي�ĵAd�4�' X4�,NH�C�b��d��g0�.&d��rd�����٦Ir�,�U$F�ҥ� 3ۑ5 ����B�s�����s�R7=����no�Z�!���кR��v�L�8�wV:�.0Qj�!�3�LS(9`�YQg�HVC)�������wJUE��P4)�T�>�>�k�e�3��9�t�Љ@	���9�2|�9�ջ�|6�7ސ��b� 1�զ
�eAiJ]X��E�g��z.�<d��ރE��54'|�
�J�h<�4�=�{����ji�f_%U
���xm��	0�js���r��z1�0����	�-���Ȏտ�$�A�u��!�