��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[<.[tӒÓ��
ǣF#�w"���˩�]��<-��hojA6�yX
՚AxbK�Y#��&��m��Ƚ�����'�,5�W��۷�sM_(8�7B���B�|�܅V�Qf����N����R�\�`sewp"e7��4_���n�td��FE/��Z<k�?#JC	��RHsu�����%�5�[�'��;c�ja���&(�Q�8׻��ο�S���W��	Tv���x7/�Cx��}ڜV��L߻f_;a$b9RV- V�r���
<�����>��zE��%O�C���x�TD7ȅ��J ���C���6��+@=db��ǱN��K%Q���I�����$�Z%�yF3Kd�/��v�Lm�����UN��Ӷ/]j�/[@�v������
������	��Ť���TD�x�\!����ߕ�o?���&��a":�+�-�99N��uh�Z"��ehU�[��<�7��r\j��Mpt��!YGBb����7$`��W��TΫK(����vK����BT��MU�V�c$�b�HޣU�E��f��O�r����y��P��y)�K�Ѿ?��TS�_[�����~�10�+ƇPu�`�*�t������A����ݺ��0@v�'am����L����1��$��f���<����"cj�d��"@�큸)N�Ԛ�)��ض�[\���g֣4��JZ�>�2ўFϰm���i0�N ڵpk���uG��B �`�ӛ��N���6�c����K�����8�W�#��_(�p��_��
�r�G��*�҂����tn����&�^};g2���5�T��t|�S�S����P�d�)%�u�3=93�#��4z���[<z)=�f�<�]�s�z*�������F���DGp����x�O��]ŧ� 0��y�Y�w���S�Y��|q����}��^��ޘ�BVPP��q��J{��.rf"�o���x6� �������Q�_U� �l����a��ێƻ�f�z ������4U�k��W�T}=�y+�ً��Vm+{[I��yRο��H�3g<�)�5��e��^�#Zd��i)�]~��k k�~p�,m�q�L��`��N�v9N1��L �SX�Z�r�a���}�ɘW��"rV7_j��������{68M 
M=�O�}�])_	��@��{�F|6Q�����IIe^� �+(F������l^������C�)���엸<���V�TCؿ�*�:�}��9ߕtѮO+c��X���<�޳��瘀�(��Y��U� ���� ���$ËcZ7�uοJ����̊�����!�ԑ��S� ��NT�:��[�r�E���N�,.��3��X�vٶgv�Kp�Q�tx7�
��4�M���(�����!2�e��_�0)�.�V��앳BOV˾���l�'�FI�m�+!��t��-�N�B��n�L' �������R/����6l�3��''�kBvI3�m�!s�U���������i�#0�ۊ���/'5 ���h���)�aQU7���/ ��p��r�Z��~ĩ�۝���XDw,��p3Cj��;������������������{g)"g{`�D��&W�b1V�yy�:>���a����I�}��S���&�3s��U���lqc\�P-��')�%��!�GIy:
��l�ϝ���uQϋ�NmX��o���rl!f�aJS�Ay�R��$��Ŝ�T=T��q�z�
e�뚝�$Q�7ȭ�ve�&��qi��9�d$8�->��F�ן�f��А���E|-]��ղ�Tl��Gmf-C�b�'4�R]_�'���-=�G��/����A�h7�3 �\���t�'c������<�(%���M�.��^6�E°K�Ͽ7�-��L^�.�P�B�E�Y/�]�N��-ۣ��,(�A+�A����Q��_\��(��wΠ9��Uz^k��n�8���؁t1�N��n��{�`!fo}���|a��;x��Qa����3Ѓ�Ɂ��w��7Ø��݅�z���U��g-�ϘN;�eI	R���{c#�c/�s�a�&���P>��>����� r].��Q�r���=�,���}.)ZV�_{����	�p��K!�DN٩҆�a�'��v�Z ��������!�2�\(؋H;l1q�.�+���%~DC?*#\���s ��*��|}��h&�'��l'-n�4/c�$���M�"�=����ڝ��ڞa�e�1�M�q�>OK��n4�v��K�NxKgo�2�����v/����ӌ��i�~�
�;0K������jlm>����}F^��s�]r�8LY��?���6,�2��a�v'�K1i����dPAW���������E�8͸��`�������c��k	��>��������Y���&mr�bO���@��e��w��z|Von0[G�p���w,�a�74u5D��0��k��O�/�S�3|�p���7��5o7��x�Q����*e2?�S��M�����;�C�ͺbc��������$c4M>��o��)T��a�#V�sw&��c�O���q�����瘨���p���.N�z�F^��7�K,�6R6���j?ڈ����۲w+��!,Li����P�����Ls�u�	h|B*�2��� Ll�uG}vR�ϩ���M�B�q�~�0��l��2#u6���À�}B���P��	��9j:
p�I �f1�
�SR���,-�@�%��*E�W��' �u�M�aB����!�ѣ�(����}��.�_k��G�H�xy_�6�E���!g���&f��-F�܎�������Javr��"Y~�x�szM�>R)�fX.l��{5eU�Z���`U���,[&�x^��!\{�,?�Y��v�}����u�5s���G;$FJ��;���S�����ܘм�}Jxy��׿i��9z
P��iq�Ch���NS�����ӀWa;���W������9�;���|w ��E�l���o+��Չ,�?��G�Ch
�����ߟ@�W�S�Q�$H|a�=τd�u�
�Z�\�7����<����/{(ahC�SL֜3�0�2�Ƌ�H����x�%gR�R��ź��pN��_�C��ȰU�����Ĺ,���R��J��b+��߉F���������AX7�ĨS;D�A� �:���ik
m�[hwA�d�G	
ՙ������G2�Չi�u	�IU���}���X{�Ǫ�$F��3n��<��>��M�T��G;�iF�
i�`:���$�o�'�#B&��q�rsJ�S&ܚ�'��wZ��q���=���E|`*���e7��̺!��y�Z�f�\�w(�G�֣ :c��EB�;���̤s`'}���P>��'h��9Y�@Tj"ZXډ�d�N��+T��
���ӥX["Tm�K��'�+����cÙSh#e�����ʏEQ*.؜ IØg� �8�c�Φ���Ev=q\l�W��:��׻p?9�Rρt�1ym��)�D��[y��,O��I�J�\�P(<�'��w3����B�/�C���b��h�.��[5Zߘ�ǟW�0e5O� ��_wӉ~�%0 T��pɑ�E��*��ڏ�9�1�O1@|j�^�5�J�̐�g�?(��c]f����ɞ��=y���B2�U�*Y�>9�6�9N[l<%U��	:-�\�K|�i��ȳ	��\��۾�-5�������k��sl����/�����l��Kv�x��|��.e�P�����!�c�~E�()Pۀ=������3�N��Cg��n��GT��	)9>��<���6ml��I-"��{N�Eec� ެb�|1�����eJKk�avYc��km����*4�p,�0��ֺ�"��a���Ij7|���h'����k3M9U�S��i�fF�&�/H��l�I-�W��"�y  ǧ,��wV��+��0T�GZa5#�zd7������c�\Ɔ��M�<�0�[y�4�(�S�j�~w��sS]�D����-�����r%!6�1�0�.;�a�31wr6�Ǡ�k�]9�|m��tS���B`��N�����A��d9��h�(r��ek���,���q��fޞ.s�� �2l�Bm��s6�ߢ% l�z}H�(���V�4ۺ��Au�1���R�4(�PXe�z�.�����}�Uxo�'���׎�8�1U�G�w��L���Н��*��}�t�دy�=F���A�u�s:����}��|���I?_�L/3��$x+�u�#:���!Zh��n����HnK\��m��:�&xL�y�2�â�4�rѽ5f,8�=��r��%��{(�����0#�ul^Ʊոp�
��2>��9�*��ݣ���j�!���9�&��@����P�e��mOh�����p�I�?�&e܃HM���3�7E�S�����Y�9�NZC�Pa�bx��C���Dx�7��b��t$.�������A�Y�'h�:߄��l����Ã�Ø��O�=K0;?]��ڎP�����H�R���j|:���cE.�em�������D>�q�]M�o'���9ܝN�����*r� V"�(n��W�jxϛ��D��������[�q9s��g�6٣���SR�?���JR�[�vJ��f�Q���a�l8��
�d T5Q�z,���l��&^$��ٓ�ȼ!����o���k1R�/t������M*/�MO0K�-�^�n��1�G����c�'Y�!7IƢAM%�f3��9X�Oh������PqX��N��z����f�d0~Y��u=��nV7�$�aM���{�Ĥ�a��Z��̂���1tm	uw��/�0����# q�j�·S�Ŕ/��8g ��Eb
�EX�D8/�':xFC���B�h�<Wm��#�q�`��~hZ�X� 6�ćJ���)%�/$+�4�]=����2B�!���Z����+b���<RO��B�S~�����7į�Y�`?�]�'��c��||L��F (V�_|$�75��^��wj��lZW�.43@�ا�t�Z���֚����)��TPL�?��b�2�;�Ck�B$ʁ�Ga����+��G{�j#�IӃ���QDZ1K�{c*��PSAu8�c�	r�����/�XI�&�����L�$��ӳ���7׽������흕V�,�*����W���L��.�6z_Y����K�_։n+��tĬ�n\��Be�4w7(�rZ���D����YE�!5�s9e�Ư-�C �.�����fBc�M�Ɖ��a���a�>,�@ձ}��|�П ��T�/����/��Cr���jhƧ�r"]W���u�s�P�+ۇC�������e�}K����#O-�б��;�{(��8/c��;;�<2MI��.�����.51!�'ַ#�9𫩁�N��*��˹�Y�lD�a8L�1S�u����\��*�� �` ����oC�E5��[�:F.����@��I�����&��J�~�mK��9mzdH�3斘rK<�-t�p͟}�i����U��m>Y��!����ѝ�|s*MB�\@�����b����jH���� K~�Υ|D\��33��	ZL%{s@;5���+�&�C�����=�<��w�r�u{�ll���AيJ�V�M�'J�k��N�a�]�U�"��.�a�?����;��E���Ω���l��d*,���$X2$��x���{M
���T%J��Y�T��Ix���#2r��&6 �QbY3�}|��z��M����
�V�c�K��Q�0��B��-K���ў+�����2���������E�Z�}��+ǇټUOc�*��#(�- R�ߡ*E/<Sڍ�`�
�%EIk��X�M�F 3��%>���х��E,e���u]�5�r��c�Ra�G�Y�+s�<%�*;At��}y����ܣ�+��Y��p�Nw�(�%�W,{eJ�s��F��I�?�bzx|�jpc�<�n
K��8�>�7;�r��(��=@q��]p����H�Qm�x.��ݳ����e|NS���\�z����Hϋ�k�k�����b�x���*�p7���2�zڟ�>�R
I�Q)0EO³���g�ج���%y���!�W�<ӂ�	O�*���`���+�9���,'TB_mI���4��Qy׽�� sH���(T�?!z:fY�O,C��f���]�T�2c,,�x"��%�����$Pi�ō����xo���e#ԏ:O�GW�Q��ˠ�aa�	��6������(��=wA������R�F�p8�yʔ�#j; ����\�:5E
�>M���Z����{P��������Խ>6$��|�'q{��H/;(v��<	�\��-�Y9
o��â��"	jj��1�7Ȫ�b�:;�Ʊă���v�a���B�"�y��jm�qy�x����"W���u�Z�C��!!����?����J�Ԋ�=�<'�.�Z�@�������] eh��t/E�̞k�B'�n��t��]O:�x������vlm?i4���l�:�j
�S|��r:c@D;S`�z�b&���-�0�;����F�㑉�mc+�쌘�4cNq���uD�5K�v��ڻ�r��ܱ%�Z�����6�)����JQ��q#��X�p@�]����ln;5,CQ�oo D1�S��D�=��=��VM���꧄�td���������xtfg�?IPW\F��@�Wz?���rS�/�r��^��o(�q�V�q�=2����f�$(�O�tPթ�����Շ���%aż\�'�I�3���O<��_J��C'!�!��et�M.�`:��Q�.�~;s����H��R#����s�&n)�-��Czu��X��L|��.�b����$�A���|���;�%=�}�W��%�\��Ş��(+��F�_���*2R����L�#��Z]��4�^�;���㯦��X�\y@q�-���K�62�����vЊ����V��fy���qQc��|h2ފ��LCM$�s�t��2�x�Ro��TcG�]^���:[�Xgs�[wmj�4y�p�I��M������SuD�N$c,Zg�)ɝ�A!�gb�+un�
ǺJL+�M&�0����ϔ�{�ŌlIJ���n�a'�k�c��~n����^w�o�$��1l��*\��1�����i�*kSX���d�Ңx,���U�J�L��U�rDx�d���0����P��@�r�+��3PK�쮀���r�}�C��A*3�7�ana#�s�$�`**��L��1�Z�$R���xb�����4j����<��h��u�g}'��|fv/�X�/l��2y�� �u�x1��|Ydt��X;���~Fu���_���BǞ�zD�qJɹ��6�9A-����c!#��trn�v���LX_PZ�8<V�1�ҿ�t�l[S\��v;�O��֐paw8�=nH�"�:K�9�%�`��\�t��|�����N���͖�EFc�QH	��d߂�n�Bl>CI���O�	���a!t���v6�Q���y8"Ѥ����������]��*�E�M�MBB����?�0���\�{�2��X�x���	��j�qy�}�1���2&z���B4c|�����;��ə
��9�ؽ�̐�����6���3�&E�=a_�(�s��yG��"8�uF�~֑L�i$z!�㼥LX���%�@eĕ� ����,� {T�b�*���ʴ��f�$Y1��|K�wO,�gmu�D�*ΈXEʮ�a���o��R>�lEJY4���O�ͯ��e���2w߂C�f�6��,a��EŚ�kv��Rs8hH�;~���D�=�:[D��:R�Ԣ���-�*A2�,F��h;�>.���NpcI�-�m-���ȟZi�.w�+�\K2Ц%�4�|�%�)La�
yN4\��NE�qTF�mIm˕!�_mH��rG�_د���#�hM�2��jx����>-*݈���	,�f��.��V`���03\�����Bm�)7��zǟ���[J�V}\���Q��O"X& eS_������ŨϘ�0I��d~Ab.b���աW��ی������]L�5�b��s}��oQ~~7߸`$JA�	E0��F�m�D+5�c�`6�!y�~  �5���4{��T#[0��V F4��H��OΝ,�%�#�]]�񭈞�x�F�E���j�\��Û��ٰ�%m��%3�϶�:���w%C�Gx4@�m2�%�|Щ�~�3ĭ��vG�i�4
+�ɚ�q�����>μ>vc����e��,�*#B��d`���m5|��k��/��7e�E�TE�\�9@�� f�@m���SH�Q���
6���$�N��@z#WJ�z�!`���3yUǘ��p㴾)3ӭ�Ԋ� s�n�'��'"3%�!�`j�$s��� I�s�V}I-̒b�1˶O�I�ٚ�[�p��B(��� &�c�1��/rY^nͳ5�x����a�]J���0���}kSA��N�`���������G������"Ԍ��(�on�'�لq��]��YY��8h�PR�q�b����6����G�ȪN��)���>���Z�T~��O�)"��!�Վ�)o���5��"�8�ll3=9��t�|W;a�mm4E(~��� �0N�JZk�� #WYgy���H#3�OV�`cY"��}�h�AkՀM���vv��#�6fXK��-���,p(���>��E���h�����o7�gN(�b��{I	���ev4z���c�$�,bR.<� �$��/�B��,���@�`ߊ�wncԢ��fL٭�a<G�t ��IQ��7�K���I��&���$ty�_��M�_Q�*�4`z-){���)�b`�L>�<����I^Q4u�N	�.�K���˺o��$��Ŀ�x�f��g������i�}tt�D*��[�||�������PM��A��q� ��,��#:�cI)w%-�+��W�<�$4L�����b���}W;�U��s�,�p�IU����%�B	�sNIb�;H�)������^t5�C1RОbRuF�����47��9���z6�ڀ:-T���	��k�t�+>�Ċ�m)�I��1h�>�T<]�H���I�;��Ҁ{I=�o� ��R#]���f֞�1eh����nLr-�7w8P|��":��(8�7l 1.G��-�\]Q@�r\��H;�׼��SP��|���	���3�0e�[������*����4��l�Z�'Y���F��\
6�&�/T�0!W����e��ݕQ��3q�"Z?l��񯃛oU�:�\[n��m���8�ۯ���*{(cd���B��?<�h ��|�d��.��D0� q�eB�H��P�@D��7M nAS�w��2��(XʧBf�4O0�q:�VA�Zi��®"%�sSp\��9�^�ջ��\?c�س�o����e �}�\�)C�b�@���$&��/HH1R@�U�?,iN�y*yA�R�o�k�^h�c���=^�d��K���o&��U�`&�p�څ�v�1�z�����}#�8�G��r���ѫ�)��z��Z(o�f��^��ϰU�\�����D�v���w�-G�J�=�r�-?�Q��_�j{l<h�9:Vk�B���zu���1�b#��o5w��)�?��
�q$�wOf���5�=T�&�M���N�廘�� ���X���k�Q��o��E i5E��O���ӛ���h����\j��BJqm��m��]/U�-K�9h\Iwl1p3h�w�5��*� K�dM�><�!�8�X�KFD2-<���À�רV_��n�`��8*�.�HpQ]��z�a7Cծn�ٰͯ����n�J�9̹�������<<�����/�"����*��b�?�W�B�!����kwW��B�"�%y�fi��u��%8s[�����PK��U{��!�l(Aë*c�]�F}�qU* �7�4�l�9�DG���8�i�;�6C�io9#f�����-���\-�*^I���D����_'���=gל��	�]�f�z \�B,_���	^"_t53$�޷Z]vaV�D$�9���_���7��|������3i	����S�r�ޜFYICղG|=�*aP >�D:��� ��_Q��{����n��}��g�2����t�VZ��l`�'�:� �ebh�!AƖB��ՙJ+��i�%����䯧�3LB+q�M����������_e����[�gõ���<��	P0