��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c�{���	��%Ӽg0	F&;me@)]Se�^�	$�%�v$J<��bݠlU�e�RJ5$щk�z�l����V��9�B����i��΋������m���������t�v	<?o�y\F�n g�)�V*���|*��j�J,�ä4�E1CTq��b�k{�u���,	l���'��>y�]8jJ6���l!���m�8D��)����t���q�����H_ka\�琔�>|l� bU��bs��y�֧H��u�Q�E�@��?��3�|���xB;Ԗl[���)=O��qp������ySr�-�Щ s�8��� H�;����d��(]���m�S�C7�:6-�b����p��˪�S�+Ռ��[���HQ�U�a;
�^��f>�U T=J0��e-��� ���̎��;c,����|h�����D�J�F�+��&ME�$N��@�D�w�'�!O�f#�FU�)s#��HK��W~J�\�c0�P~h{d�T��|in~X1W�Y%"ն���� ���B�~g�|����k�'�*����T}��H��#u������*u2��{�&�`�VZ�'j\r�x�h��k���7�w���/x�p^��)�����B
bZR�gf���f
mT�������.��N����%hO��5I��x�T[}�Tⲭ����{`�{�)��]o�h�}|��wE�[:5������c
l�����5,���[���]��\ Z�
�X��ڏ5=��4aK�E\L���S� ����ش9�q�QŪư	��v��Z�=�m������z uƭ����E�Z#�:`�v��e����Ǩ�����m��.ԛ�#N�[�i��؛��=4νЪ�q��H XW����)�
���CCS����9��j���E��!�/ן\��0,��ck}q����ϴ~ ��A&��R~ 7�m/�d7r�p�@��1�j��rf�E,`S$��Tt\. H7��D�h�k���#k"���>	�c���aG�4���4�����ק�K�(Y��3�_6!�&���4u��[�-�S�e�Lt�ܴ3��X���p�3�!8��s�˥��+��}�b��vmq��/٫����΍�ӶPĚ�gl���~M�Ҫ�W�;�>+ ��ǵJr��¼E{;�!��M��q����D-Q3�X)K�'jn>z�>�=�P�Y!P����Oz���JY[d�-uX�~�����$���0`q'��G�����[�Cq�T�S�8�.0�3��J����1��:�����Y�k��i�d6�5�����'�'���:���S�I�X��眔�(��T�����᱕ �e���Ρ/T�Am�+�e6u�X���r����~��آ�`ŕ�Kp�kq<r��	�	�U���d�@��-���*kA��Y�3ճ��i�&��{�d.�t)W��I��^9�'UQ�t	�Ww���}W�}Y�)K������V�B�{�?�l)�C��~�5��ؑd e�k�+&fP���Kj�̓A��K����
�aH�����q�5#�!��a��>��|���_��g�2Iq {���)��ɟ%���+��au1#�	�IӐ�w=���o-��jE-�����zp2����������I	�>f�ufиbe�J��اc�� �S�<1���9�s�Ͼ�6���A�5��/;�vh����bT��,��TXC�y-8
�kN"�5m���%[Zø�M|��j�y����Й�q�����x�Aa���7���soV�1����v����@���R zȓ.9I�q���EqڈC;<�6�������h�{�إ�E-$.��M���W~���v4��E��me�~,�%ʅ��O>����9:Z��8X0׬>Khw~5c��j��RJΙw����-���H��Kd7�#��7W��-�,�0��9lhO��X�����d�F�o�e	n��g�faa�C�r(��**֝�<����9;�k��=��zm �	��=A6F�.;j�t����%�|���TS�JS:��sk�F�q܏h�9�\q���Ÿ[���0�"W��R�+7�@I.�7��-0&!`Sn/��P�1d���N
�Mi�%^I�TN���ۛ=�Zio��f�#�l�+h;���V�}ʫ0�j�9� �Q�KB���g�h��
�g��� ��)_Ր>5e/2�n�}�
���h��iѬX3������4IŌTǔ�B���&�U�G
y�6i����Շ-�Cp�N��Ja<V<��#�����Kk���T���{�Y�\��bT�k��,9�~�u�����eZ���Y/���zBB���v��Ir��4�><'8��{��#	;8�a��z46S/'�c7k�*_.о�(�~��l����Ɍ�E+N�>K�"�A,(o�lf4u��_*(l柹�|�6� A�hPVtA1Ǚg,��{���, e3v�|+H��ޫ�W��n�K�P�7�7���ĵ�w�L}��l<��F����2��KI>�̜D�7x�3�\���p����9���!�8�ݍ���;��X/��!�&������b���z�oԟ���^Pr���%I-�3,�8Q��OX�t��?�����cqb���=��Vµ߉���z��Y"'<2�졮�`LY��)��WM������\�\E-����ʰ��j�A�4�::���ր��s?˩����(�ި�=8�j��P��"�c)�r���#Q�g�2F�����ʕ���soT2��n���h�q��� �)o{�E@7����Ѯ��C�`P�p���]H�e�J������aQ��W���[K>N�k3��_ȵ�o�^�uW���}�\	s���Q���Î�r�zH?閤��Ta�;{��^�"�h���AjLC����=�V�[?���i.A>��i+gǋ��J>A%0F�&��~��+��U�jf�Q`���[�����]{����S�=�8���4	\Y�Y�/F�
k�DB�q9�>���>��V�c�By*rnD����H�]{�U֫'��]�������sDVe�Cn�H�eR�D�Z2��ʭ/�a�ȕ�j.�mX��y���lP�~��[��W��|�ϊ��B3՜��.�l����ޝKSL#�ZL�
k�D������-�odƽ�(u(m��MĜ���*S�(ut�8���R��~RK.`��L�z�.۬~ӗ�T����|0$�3_�?��C���.�n"��~���̳o*f��	�<ل�HǸy�9��ǌ��Ɉp�2�2�yY϶�� �ÔCGݷ�(�X(x�D
ڡ�@��0�_�(n##�Cz&�en�v'�GW��L&���_%#��53S��CBS���R�ͪ|�L��G2)`6�Ca���Y�K�z��1�.��1c�fs�h�o9����ǹ�Y?�sZ�p�g�$�A@2�%���\�U�m=��-�xuc�'�j�5��Ŀ�K���Y�2hSD��#�׻ hv[����ͫs�>��ѷe9���R��^��w6V��?Ԝ'�P_�C�C?����Yv���A!�	�ڑ��-��&A��AT�ʳ��:SM�箟��-܀&M�u8a��!P��������nK�V�&��f���A�t"�M���*�'7�7+�^_O�FQR��T(؄y}i1i4�ـߋz���ce��QE*�� 
[.r�("&ׯ͍S�N�M���Tݛ}�w�3�ctu�*������H.6�h6��0I�MiV�p.<���j��h�*r�vN�e������"����@d8|/��J���x���j�r�#Ha,F/Z����c��P'���Pm*�'`A����C��)�-B3��ܭD�0"�t��.�F<��o��ݜ��~�-��!< �8��X��RMۢr 6yF�
�
]��݉��闺Is#���鸎y�ze�T��[�������_9ߋ�W�>+�VOl2z�}^Ďv�]�n��&��4��W/'@�Kd3[�굒��2�XU����.�5�N�OS0��Sɀ����M�����;rf���ϵ;�M�k�wݮ녽��B_�Gy	�H_YH����va!��e�8`g��{S�2ݬ?)��x��!��0�N��.����e�c��'����Ϛ��PT�<���|j��s��ߵW(������nh�e��"����^i2F�hq�]xـ2��ݷ�>ɗw7���O���$>ʒt}���=DN�$��Mu\�!��Q�5������i�-H��;���.�g���%N7+�z��T����'ո/u"�1�+���]�e�!��h<xL�/�1o̒N���qz�r�@�S���UvD�U�f�ˎn��%�6J_��ެ�Nl��#�R\�d#�˂o�>�$�o�5̇:���g
�>ƫk������W"Ƒ�"��`�*5��k�}#\{�gr[{���P�7q-�	��6�@H����2x�%j�˿�ю��c��c�wk�>�	,����`�7�%���j���e�x}��>Δ1�4�m������>�s~ّ��݄+�چ�X��G�8d���v����ٴ�[���Ot�
�]+GB�6=�I�f7�!ފ�u���~�L�DШ6 O��QC����A�[�u�ȃRTF o��&;��VR��,�C����lJ')=%��G�5=�ܩʳ�~�cR��bh^c���W��yqB���Eؑ5�~!�tS2-� ��Ft25��v��Uy��Ϥ�wG�T�m5�fb�;7��z��w��5_��@��P�g{� �����G�*:;����j�r,Vg�==���輿tg�ȧ�l.ʷq�@�a�,ū�s۬'�d���#��$����|$}��x�1�=�FP��Z����K6
SDNP���t쬵�m�WW"q��e�X��>��w�� ਗ਼�k������^t���ߠ�=����+��
7;�ԼTR^O7's9@���,�P�����^�XΆ�k���h�(�oꑔ �Ō��s�7����Z2c�2���*LS�o.��Dw����0�Gڜ��tJg��-�=��ݵE�`�<�-�q,��$���=(4v�ȁHU.