��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cЌE���Mmc}A��J���[�UN�>��f���X�y-���9dW�j���ש�3�{���NB1�{����^V�8}���z?<.�Pr|��4���o�E��ZPm��@�}����\��d@s#`�#�-]�m��V� �H�fP�j�e2q�2���@!]~J�z������M�2w�����WP��Q;9��ODߤKW'�{7bl4=�K�(��XzK��S(`f����|�'�CH�����72��!���01*���w��Bg�Eo�x��$�
mJ)ͬ�����4�2�z����$���^�b��6\�Q��`$]�42�U�EE鱘!�d0g�ܻ|�-��P}(�[��=ڑ�161��o0��{��\
�����2�M3���;a>T>*\%e�R�F#�� 2k����� �6�uP�����4���u����c��!��j�J�ݪd�JDd��j�h
�w�����Cԇp{��3���L�,��C"�����хa�(cv���u�}��a"�P[:d�h�.
��-�0�cZ��d#��֨�x�2�,rK���=�D�6i>�U>妥�&]nS˄��� H�rW��ȴ.n���kW3��mP���䲾����a
�t��?��֒�ƺ�� Ik!EMO@�-�X�����W�a��������y��O�h��X�~n#��e�!��������)4�T[����Uu�Sv?�E��9I
z�rr�����>�J�a����'�HJ�У+[�9���)��Y�`�7���]�����A7�b%jZ����b��bQ����66�k���Ro��� ��%*
���ul/��Y����e6Y0��=�#r���ul�{#IWDjE�"�D;�U�OYj
#��"P�b�s�bj�����2�9{}��~���k�������d��}� �G:�l��z���t:0�k����/k��L�ً�+�.�U��c�B������:@5��x2J�=&�=LWCѰz�Z���h�²NY_���,����h�2P٥
{/�� ��>�F%X�� �@���q�6D0���%@�CR�Je�3��ć���NRH�!u&7�%�В�I�1咰�,���G���Ղ�N8���8z��-6[�e�?�@��Ԅ�ݼv�o��#�zM�24C��S�\I8τ�e�RH��%E�Z�hd�+��3(f��ήbY�l[;C�k���&��ս�g"a~l=�����������:�Y�.p��O����5!�DYg����Äb�6(|\S��r=���ʎ�g��:��Iy�ډ�-�8&$�E��F ���r��lGD�)?�D���m� �/���LCԢ.�e2��~sf|�p�@�m_H�>#���3c��H��b���$���G!�N��UD�9�_�J���� �)���0{]Mrウ��I�'v�dra�wE��C=
��C�m`���K�"�+U�N�i��M_}��MZN���z@��>cm�Z� �3��֌)it;lƘ����k9Q6$n������%N���,�S%��N4RHes޽��S)}1.w���u[č�K��*���.'n�a�&�,�T"� �I�D�8N�S)�x 	�d�;޻��G)j��D����*	��@Mp�sy ��<�mm���#����J�aU!�pmm��7�.�`	OI�{T���9N%�(��������D��=1��-����IF��˽ЗO��JkGC�/9�̺�E� �j��ܠ]�x�֒2���m��2CBB�jN6؇����̠��x�FS���-7V�����l�!�z3l���T�L ��:��ǣn�Eu�t���	����@���~��j�C!IBM�LM�kg)q~ >�~^�����,���4�,n�y�$�bd�T�,y5ҥ����,8xnC�*j#Q�D,0��(��.F�v�<U6j�����8��ԙ�뉈˹��2����ēw5����c;V�2�zJ�1-�4-��"�����,���e�j.�VpJ/�p�0�`U��Z�C��=-�w���o�[>��o.���!�Τ6	��v�Z� I`)8���y�e$�����E�=�t٫��;N1�0&G�����"�'�o��p9K�b=�j��ii�L�XZ�7UM&����,M��0�J���ȡ)}�����WI�|���O��E`�