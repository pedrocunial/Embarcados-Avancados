��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c��5�h�:�**$�'L'9J�k��DB���a���;Qa�P@"��՚OG�I��U.�?�R�ð��y��j��GIK����w��.6��
]��9����޳pI�@
������O9?�C6�`����i��n�Eˑ�Y5怅Z���X���0���$�聾���B��h���j253C�e�]}c����(��EF����(��G��,oO��7�d8��W�1�a?��w�]�\e�V��ͧ��m��X����r���i.�ާa���������O�n	�c�G_�����j�??��x�IY�0x�<��_v4���]Y�G��7���R#���7�6˟�D�	�e�B�ܯ�ٲ����(3�'���T��HH��$kM��5f?i�������7��97���(̱��gWp�+�{�;�*l�s`~�m�,aA�x���<5�����h�(!�<�v+�E�Y�E`A���t���hZ˲�	ֺ�O�d, ��?Bx��5��ؽ��g%��K���Y�>ƓG�������*��k��yj�(���F�M)�Oh��I:L����- �u<��u�3��p�r=�t�JG�B�E�2[�tF_�IMA�ɦ��)��\���ԡ�_�a��~��hL�{���+���A!Ε�C�*�R�ؒI�uA�y�h�D<W�e�Ȩ���C'��Q=��d�1ʺA;� fq����;*�/�p��~��*�dҵU�+�`�bwQ��/�\��y�3N�\E�%��Aֈb%���*��'fl��c�O�4[|O��2�^Z��6��9�M#V�þw�Bٯ�S�U��"�o���ߍ���l׌=b)��4��y%4���|�) Xdy�1�Q��àa��\��k��io��u��(�޿�x�����w�P$��j��yT���j��%( ���n���ϭצ�Hsq0�b�9�ք�F���Y�a�ji�~�Yǘ��t /�_8�֌�����G����P�B��ڼ��\+�t�w(v��-(k&�4Ud���n����8e��>��|_k�[�v�4����h�ț	�-�q+(a-:ߤ�5�̭U��m�G>c���ۨ~:�7oؖ���E�l�����F3�G��;�I)���gn�a��(���a"p��A��h�sЇ�h���gp>�эTk�km^�F{-��.���ֲm���4_\�	�� �v�%�rK6�ӕ��&f�.�E��w��$�s�-�-d��Xv8��_%>ؤ]j���bHo^Z��H�mZ��Şz���*���>I�^���34a�_MQYW��4ǲ>�ߪ�k�Z$���dñ��m�%�D�'��A�J���qp�0>�|�(��'����ƥ�ӈ��������n���[ �#��#a�L�O���B.���)��D&B�I���,T"y��M��`�0�U��ɥ�罩Ld�UPj�tE#���Yw��:Q��.Ｌۿ�o)�6m��B��KnM2(���w4�Kͤ�	0۳�
�s�8�صl&=1�)h矸����=�;�+�m���O«��Ǜ��U�3bt�0{�ȗ�t�GSD�M�"��{�e���DX�(Zx�ķ~��@:MWE�CG�U2�x���I~ ���(����)�ZW����6��������'�1�b�l��&)c<�^+�/�-�u-
|�~�����/͊�ι4.6+�cB��2�BufE��9�Ry����eմ���Wd�9^DI!&L�E]��bah�9�����=@bE��'�����}M���X{��0@�Q)��Z�Y���eer7G�/I��TK�l�k╰�ә�l���6�NԂ 8�1(;�6VKm���˒RsR���ga���
�����	���S��ȹ|@��`����>N�!�L/v~��U�wiR�'� �6��EĄʜ��r>W˺��X���熳����ɛI�n�+�3?���I��
3��楫m���Y�*��2a��8j�V!��κ�,d���r�Z��`Q�ڿ%!���u<����Y�ơ�6D�hh%��Sjƪ��<��ܪ!2WC��$i[Ù�y���:��O~�ˆ�c��K���V���X� �:��͛ɟ����. �زFW�F��.!���V�Vxs�tW�Ii#�z�[?�`���)01���P�jB#5�t�Qn잋���kr,��S>��ɺ�h=̐���� �CC���G�a� ����ZQH�t>
�CI"��Ͷ��f�~�A�)!�X�l#ֳo�/�!ݾl`p<b�u�8~b�Gt�#�{�Gv`���:((�km��������Bf���Ea�KʰuF��ESr�ŷ�I{ŲZ�xo<���\H�>ø�Dd�:x�^	�W�t� ��t��R����7�%Q=�퓞t'B��cP�0j�c4��M@X�+��'���6����]�3iwm(�\��k4����Υ����i[˷ye�&ʉ*P9l��Q��)r�\�u�!nhq��ʲd$p(hɠ�.1��W��k]�U6O�Sm0L��1���7���`�r}�繨�{� I��������0���o�`L��4�ܰ��K�j�?ï���+q��nV$$�����(`k~U�l����I�O�!��^�*� ~-��\����0�o��ߑݓ:�oh;�����sP ć.Νg���;Y��q�ǃM�Ja�݉JG�S�,�pd���,b%\^��tlfB`|"L�.e�NU�sS@�Â��0/��f��s�r'�]�����CN���,����\3d��"���a��#�a����A%�C�	�`c�G�틓���Gϛ?�X�I���#���P�C�|�6z�1�в��hzٿ�p7�u�݇_,��bߖ��S���PV+�0Ṇ�����Z�F+~(L��@�1(\�`\�M���)`]o�0s�{�ռT��5Z}��یCQ6���{mf�����(��n�Y��DM(���;*���ZN��3=�~�Jh�{���9! �n� [��4�Q�w*וk��d7|���:�~��J�SZޱW�tk�QfÕ���7{;:�
)G�>�v<N����C\yv�vP��gj�v,N�3�ң�D�����y.vgBⷷF�xr!� ��]3nz�b�k�巟g>��&�� �{����8ML�=,�f!�IzYC$�+�^kr�&��+��G�`%�<g��H.�_���0d_�(�F2��!�QhyN{���eYtp5��c�u`x#�V��H"���`���+� i�lX�Ѫu����V�k$kL�O+�a��aҷF�Aڒ_������G��n��:;Q��~yF<<-1���Q�LިҢ�Y��cJ��yH��X(��l*�a�U��$=4�ob�c S�*e�Z�:\O76�AXӂ�S%�3M�`s�w��l[`���/4F�=`HӤ����<N�;b��_=�|���>a�:�E�����*?�P��e��LRB�i���! �B��'��&HK�(����zm�|Z��?�X���!ۃ���њ	���+C��˘�!8EV
�ɳ� %��w�DQ��ԅ^%v�
�@���D��l���j���*D���jO7x0�2nCYvSX��Ɍ�R�i�pV�f*:�f-yZ���@�$�7'��4)�`�ضM�Ϥ���0sq�w�T#�^=F	�J��Mg8443���S��qc�&�$��1�-)Y����<�^Q�4,���ˉqi<�G8�nH����r�����'uՐ�5��"���=�Sꔙ���0�\Sȶ�U��fJ?j(�rl�|�z4nrs�S���=��d�;�j��v���4�ͼ��v>�\ަ]<��W�Բ(�{]�i�k�Z֟�d�[Ђ��N(��\�o:�nS�ڹ���d:n�����OH��X�6���l�[� ��DJ���0<Rb�d�����Uy�QI@�y3�����s�]��/�{'Q- :�a�n�Fi��ɰ�Fy���O�"�"�l����y�Nl��M�u�f_C��oCH+��]��S*uO#�g�:J���U��!,�߳z���Β(�Bx�Ȝ{b��?��I�}S�3�����f��Hi��*��b-�F��ed�B�����6X�1*��"�����|:�Z�D=�q�JP����Z��Ca��]LnM2=J�����5bF��W�%����NnB&aO����Uצ�E"�V+��)x�Ðj�������@H��Te��Y�����~s�{iLh�&+��{U��ŞCν�AԌ�?��|�����|�ƫ'�*�H�m8	р��d�^v�4��������vs�$�k! �X '���
HƆx��I�(��M@h�7CP(�U��Z�軧&Ju��P�M-�q�>f}U�����u�B�֋]�T�ϴI��A�}�)��z�����i˻y=*���k��%�e�6z��]���%f ���88!{<@a���my2�kE��I�;f����=kj_�5zS2���8�����6���O�*{Ϥ]�gG����2C�F@�c[:��^�tIǨN�:�㙗��$��flCVԖ纺.���f߯���yK�8���w�����,���oW/��lُ�g�3j��,�������i�u�||Y����V�<g�0�� ���j���%1!��]ड�sP?�E@��-���%چ�-�LY �|��{���?M�s�Q�ڿ	yV� 6h�)��,K����,5��V3������]=Rn�,�4�40�P�J��b�I���4��4���.R ���ia@�����:��G���W�Am������uԀ�dx���, %�5����G7>���j�`л�y����
��� ���{��'�?���X�\w���"���3T�Վ���?5��R�D��J*��RH�ý��%�.A�!_Okq�V��F�5BO��^��[�p�J#f�y��5 ��COOi�n��-~I�d�z���Pa� i���IC���ӆ٢$v�x@�ڻbZX�I@MPʮ��U'0&�LbQ�:ַ�9��Q��4�O��m���n=8�����&B�6͟|���^�����:����J���6Z�[.@�E�n�-����y����O��y�
����L(���;$p�3��՚�ӻ���B�o�_��*�z�mz>���gl��r���S�Q&�H��I	� �L$�����Gh�¥z��)���k��z���X�=��M�N�݁l�iQ�8ν"�{&\Q���%�!4ê�)��s�����j���O��D�nj 5���NS;�e��S�U�ѐF�^��l���AҖ1���93��]e�$`vI��g��y����aY�5/x�--:6gE�x�}
�A]:hpـ��U�QAX��I�c���:z<Xl}�U�iK繵#ѵ�����9�%�om�i��ș���"�\(,���dS};��ϐ�-\��xx���3Ʌ��&�K��!D��a0���v>�-������m�w�:��3�2.�._6���e�i94��Ԫ���sX}�u���*��s����/��c<�{��L�c��?JN��@���a����?�R��Dw0��Y�������ٻ���.b��eG��RYHW��v3O}���*��߽�Y��|��o㙾k�}���:k��k�}/}��]�C�Bn,Y���ΐ:r�oq�{sH��]R�|Ԑ�K8��z��ٷ�M}�7�n���@�T0Cהer��u���̳���-�ܶ������x��� ��]`m�K�G+�Xp���W���V��,!�,ӌ:�����;�GH+��l{ ��[���G$jF�x�ۋSc��Aͷ����	���uj9�������uu]�7�	b��ݳ��E<����h�4������GI`;<m������Ϸ��&]_�3b��^2(ߎr�?+J��qF��t#W�F�h&y��t��8X�	�*3$*t��$�er�j[������9m���!�O�� �grEZ��|�ʥ���qL�*����#���GC�Z�ֈK�����S�D��%*q]���bJ�5A�wU�пu<���F�Q��әRL:�� ��an<�w�s���.H�גy�u@tp{q��qb@?_T��z��׽�dP��^����ީ8j��e3�]@�/y跋�4}�
w}�)->o�]�&)'<��6H��,PP�ɫ]��v���D*��N,Kh�"�zJ�I���u�ƥ{�FR�ؕ��>(�����	�q00�a�7������Xp�J9+�+�ް`N>q�>�T�Y|2�h�d��ȬzT����L6�:/?"��n�1�BNOKP���
�޺�m�P=�,B*C i�N{`�Kt�o\��f���"@[��Go����[�̴77�c�J��@
����\�
E,1�{��ުe�9Pߨ0���ƚ��T#pnTd��F#eY����j٪ǌ=4�?T��f�'�8g]x%H����)O��U(qJ�qqI
YH!�a���Nd�#�Wz`V�t��F��Kũ�p�H�~���b��[ 
�*3 Q���en��O�#9�:��mH�������s �B��yp��(Y�|����[ض��P�T��Kdq�,A��L~j�ws�^5���5X�ܾ���=���c�������U�����=���p���!�a�>�J��y���]`�& �fI��tm,��=���z+%f,Ii�">+������]�C����d���*P�8wZ0�qa4�k?a��]���Vg�b��*��o{S��!	�3Y�롎�����x��K���{��Ood(n�����9�qu�q;�8��GV�����W�&u&ch����C�3"x5��U�j/����􆃲}�5����&5h`�=���j�d%~K����<��$�al7����K�!\ g��-Խ֫=���ʖ��?b��	Y���q6��L30`�����i��g�� =�>��vK���Y1d&.�'�]P�?M@&x'&5���c�:���{D&<�i��>��"����}�����N�Rg��'�n��P'k�^3_�|ac��h.���ͬ`c�m��ZF����5K��`c���7�Q���av�'��ep�k�ѻ�^9De�u Zw�i��ս�����&O����W���������4��.E������U��?h�0�8���B�ӆ��F�;�<m7�Z>�R��h(9�)��^_Z�eC�K���@��<�\��S����W���u��`D&�U�C�'֘ ��ؘ �� �?�����N��j�7�|�Թ���k&�',jc��z��ݔX�FǕ	�I��WRU�S��o���79�$��-A�T��rE��}�&�r��:��S6}��f�Ew�6k����ݴ)���*֟F� 0^�<�Y���<��}c�"��&�S֛����n�×(��b[2��A��G �<z/ȑ]��?�xf��]��y��3w��u��l9Hp~����4�U��>M��|�`�޿��k��5(��iV��^�Gh��6߫h[�>7% �P_��B杔��e�%�&>}�.aIx���z+3*�ǰ���u�����	[9+Us��
��ϭ0��YMI��dL�;-W�N��5
Q�[��_��]D|�����g��:�b�/c��������Z��"�0ϵTK[��B/{A���PV�(p}�8>u��G[�¡�yG����I8Ơ	]���)�/KЕT�~�:�8ڝ T�Ꮤ4��[��UBEx�"�څy��/���W������CM��X�N�~���~Cm�9Τ>�y��j�\=D%���Lb	F�c���a�2ا֦��*g
�2�	�2e�C:�qSlH���GnyP1���1H��&g�䓂d�EEk�� �r�0*^C��y!sx����ߣ�����G�1�3$��ⱍk�@1�!�<J{B8�jcۓ���R���`��Х)���o�?��T>���9`��3~r3]�},.�X�壬o�5m��u"7�6�6��ϫ�0�І��5���c�bާ��VFQ�^p ӓy��gq�/����y����:�d�G�����t��yvߒ�{>��ۑ�8Ăa+s}Q<�J��LOj%�S��꾈��eZ�rǭ�ΕӍV�Z�l����#|�"��vF�j	�@/��R�D�R�E$x����NRj%�An� 6I�+cȪܴ�>NWvE7q�������gO�g[����K
W�-�r_��(N�R��
U���J�k����$F�t+�3���0�s�q���yD�����L��މ�m���i��� Lc�^�-D�F:yy��Q��8��ӘϞ�4hD��7�Y����'�i?xf>P�ol�+��è˻Rkl���=_&k��V�d�3�K0��`$2�,���"��<GD��M�i
��s���\�\�����2;I��=�5��Y�*s@]o㐚��(Z������lA���[��=�O����n`\fE�ϟ*=~?��2IBc�pɌ[I����
8C+�ёE%�՘��KY�E��,FD�4�W��
��[B��_�3k��C��qE�-Sm!�˷ݬ�a��OWn�?�>HL�m�^e�й5���]�P�15"�=����=*\n7�+�ȗ=�gw|,J�ƮjV�N#L]@����4�W�*3��Ջ^�c\nd<����f]"\ה��l ��
���������s�;�NW##�D��	��a�˱31�ˮ�Y铧m3IbդAԓ[�s����^uR��r�o�B�T���"�qxA�|\��,��ȶ���)�c�1{ry�TaL�[9���@�!�!������$�����+#�`9�H�~�� ����7����=�Y�Qx��M�w۠�7�����e�>ZH�	A��8Ю�Ɗ=��*��8Y�+J���$Bc'*k�6��E������4�B8���&r��F��V�otD$�>чr�k���������~"i��B:�c��ZHmp}���u�v��h/�}�����'ϭz��6Y���e��;[?[v�KG�	4��k�zl0
.ޏ��H���hW3Ы�������IVIbן�̾�w��H�/񓊙��v��>�t���_�t����P�!�рo[�aldy�%9[�i��5hTep=��¨% Fk��l5�H� <��伹
¹OJZB\p�Xq�-��İ��w�>�TnC��ǅ��<d?��E���2V�3`q���'�~�ik�>TL�Ŋ+�>���k�iU#�Q�0忟嘻�6���Ի�w����(�O@��6�Y��2^_��u����Z��#{��J2�D/��d�<���B��ŲgY�<f����6���Բe�%�r��yqT��/7�#��ms#���鎝nhr�f<+JuM<σÈ��d)QT��Wt["^�����`�$���=��衕��4J������e
�!!�[�5=!p"���u��\�̬��d�Ǆ��������h�/����E�o%.CB�������T��b��A�L�*���~���4m8	��Ct�2�ɬ�~�f2
hP�~����
���E:�܉�_�>����ڊg|s;�q�T���c���6ww0�u��RJ���Yi85��Ŧ���E�S���J��(�����kk�(ݯ}\b7��`:C �~�O��z�7��[Y�VUӿFxK(%ź�inY�M�0G�w���8��9l0��M>�'��� �g�SwF~��,x��:F޽�M��71�ܦNӗ���y_����M�պgp-A�rڟ���np�¸X�cd���Įqd����eoDKv9n�Дf��lr@jZ�?Dwl=Bn���s��B3-��<l��"r,Y��;�R����\��Ukj9��A)��g��#�|����ȩ}�2L6����"p4P����D����C��V)X�F8�iYo�G^�gQ�Z���,ɨ�QeREBt����΄}�9��@!�E�2';��~d���ڏD��W,-r�^Na�ըX�݀۽׶�m���Z���.Z1��n��2��gH,%Z.ѩ5�Ԧ �w���yo��J҅���-�Ɏ�ȁbn�P����gqRTK��_��(��g�}1��XY�D�3�Rg��M���w �j�l/Z�.������Okр~m�=�;pu��RxpkR��Ų(&5*�����93���9!B֊V�w ��1:�NN7ϭFz"