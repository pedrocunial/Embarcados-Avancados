��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c���ѢǓ2�Su���;'�����)�I��߸UY7�Ҍ
����y.��Y8ŰRF��� �LNВ9�T���ag��*���=�YY�iSjD���I�*����@�	�hm�`a�Ǥ9�]b��ͼoE"@Ő�6���ԧ>~���{�J�bR,'�Y��Ř Y�i����B�M��"�X�4o�rS��`�؁/�&PHMs�r.��H�1C^܅���Ұˉ�B!�bNa�HF�f�;���wQ��S&��L(�(Z�'L2����0dIcT^��*,g�.b��ݔ3�
A

�f��6��RVQʮ� �F��pF|7T�y�u��_(��7�0�#È~�_#��έ��aJ�9gd�w����k�y����
 e���k���8V�HqSǜ&�)U����D�1���C� :Iʌ�g��,՞�,_��C`>��1�C0l��N�M���C�[w���M�?$�H�h��/�~��pw1�,��(*֎�J�k�x�
I�%�7,�Q�*cɩ�D���a�g�o��TQ�+(�"��p������[�<����w�8��s�s�~�X��\�j�sW���	�؉lV8�hG�]��EM?�uc6�?ݯ�s�?p�R'���F�\@�y`���fs&J�H�5���4������pȆL�	3�EZ���%u�դ[F�ݾO&<g���yb�0��{��ևeu8���p�/q��Aצ�X���`�
ȴE�/�൮�6sy�_ն�����K����x����a�cݝ��&P�6;�?嚧�F��3���򐥄ra��Z�[�?�b������L ���`�%L�r� ���N^�f�a_z��C4� d��[�2����I�e��U�8�=M0A��9J��{]x�o�t�������`x��Z��Ħ��t�v#ל�u~�tN�E�G�4Ÿ����&Z@T�J���1+�'�u�<l�������~Vo����?���5�@���Yoj|֍��P�E�^�|�jsC(Y?S�����F��*��a+/h����{��b����-ߊ�L�������s�`ߚ�}�������l#N�`(�̪+���Y�IϱO�O=7g0��9���޶��F���_W���N�k5tI��~#,�t��G5j;O�Ё������-�G��7^d��&!��\[W����C�FO��y��/��n�� VǇ4�iGv>���6_G��,�|��4Jƀ�
�"f2iM�%�6�!uN%�:*���M�M�f�N�cN6ڈ4(�7i�`Rm�ˀ��/`i%��-��v�K��*��F��-�y��ֽQ�� ?3\�dI
� �jU�}��)��%��$\c�pZ��}t��n��?�;
�����^�h��ꤒ�m�Nľ�~�o��2r�xծ���|px��U?�q�S�c-C�,�[�AK_�9m
.��¿�lnD-���Ȁn�M2�K�*N��%t�Տ�_P��|�u��H��nnEf�n���D(f�劼�Ρ#=<>Z[�U ׌��)L��w	���*��eg�Z	��}V;�E��͈A��	�n�)ډ�ZA����<���W^����{V�vЌr��>�S'�cQ :�Z�����k7|�J�)�C�a������A,C�l?��s�+��|:S/m�1\}��㳶X�����F��_bml�:�5<�������t�f��<���{a�������P�#�US�-+�/����!�$@��^iŇ� �\;~�X�Q;�s�Β������\�MA��yYJ&�P|��pE4R<d#�6��(|����Q9�����(xf��u�hT�&�����7˶��؛r����]�!�
�"US)�P��X�BT�;���D�Rn�[��[-HM�XJ�ط'啬��Ƞ;߳@��X�c��s"��������P,?G�f��;�﮵�(�'���w��3���\��:�����K&�.�w���^D)�"�?y$�Ap<bd�aN��l���,ݚ1�ktjzٚsDE�4�.���m���w�*�����
N8�1�v�S�A�-��I(�8eM�
e3�!\�(�8�D�S=&��C��FD�9����h)�j���uH�����L�}Y������}]:��~���]ȓ�uZ�V��8��E� Adݬ`��5S&���Eߣb�8�e���ja�A���.�F�U�8���y��7)�T�@4�ڪ6��r���kL�~�Vg�����!���3M����d�KR���>�ˈ<"S�B�"�J��_�BV����dx+�i�%��N/(�zF2
?��p�	n࣑����rAPA}�'��d�����*�x/f�B��W;����qqg�փSf�H�!_�N�� o�6|:��BӍW���ެk@�����-�h��l?(߃�I��7���!����H�O#��{FH�݊�"�l�:T�9/"YYg%���۳�eL��n���N{?��<ќ������L���f(���)z*�������z��V�ݸ�r�j�ؓ;
�I��:`Ι糏���US��W{��I~�$�V�q�o�*�s�i(B��
���d�Q*���f��-�[%��Te����d!L��$y��F�pkw��p���K{�=�����x�(��0�' �$SV��zc����o�L���?a#h�!��6�]�Й�/ѶN�p��)t6��>����Ri!N�V�~�E�CՔ��m�B��$P�K�y��>�.蝵l�n���d�o�<=ʪ���E����|2�#'��ȭ�j���\{W�j��\�k���%y*$�z~��>�Y�	�[$��6�\���!U��d!�w�{]�?����9��Y����Jڟ�q��X��U��.��˔rS�e�x�ڞ�Xe<������
5d�d�jnv.�_�'7{�Y/��W��6.�O���1���WDzc��y{U�
�[��̃uY&�f����� ��gl���?���.�Y��k*d�gW�a+1��N�p�a���Z�x �
����}�R��˨ ���b.O5��X���-���(e�F/<a��j~g��]� D���SYs8��(�v�4ZNT:S!m��+��{c�������G';g�p���	��6��CD�h�H�R�������5����ŧnQ�}���?0���)�3�p��gěx��%%��W�V�*U=ְ�|%b~��ӭ���`��rt�@R��N��O���͒34�闃��Z�	>З$�y�/��0~��m@�fVB���f�氻;d�u� �;MPƾr(��ۘ��'��^{j8k���6ia����iyD�$�:%\��`><*���.@Ch����oH�4�4^)�J�r�s>_4	��`�BBY���>`"�;�7*�{ �ټ�� �!遬Af���?��O�d����ݯ|N΅AF��-uda+��1v�����9�'��Ieh7���i/M?��+'}�Ǟ��o(���c�͋�8��T�J�pN����(m�O�IN���uL;��6�t;���*j�db*W$ok�G����jP��e+��+]��+$�P��Fw#"ڐ��J7�#^�HK'����G�N~�!E�*I��tDq���f�#K��sa6�֛�E�Y�F.�UNø�-uPE���\��Lc+�݇2�Xŝ�������X~K�kx�yf��&h�'����d���kFmm��B����d���E#�x��@�k�R�D�7�3R��G���&����K@f�q������@>�z�HX�XmG+,�$o�q�n��`�cj��}��G�K{u0V�S�%�w�0/��v��h��қ�!����̅���� �6�R_u\�K���q��;f:up}���F#h�W������8I�Hv��3U��^�L#XX�AL�B��(����S�!Ũ͌��L�:C�1��ԉ_�(y~?DY��>W��u�����_�R��~��/J���D�Q�W�,)XX|/��b+�a��E��j��5���h�������SϰX��0c����gZB`�{���7|)X�/�O:eW�v��(��!Q���/M�q���ӶFRFj�l����I�Ç?��00syΠ�w�Zp��yM�[�i5�^M�?��LS�$T�Ѯ.I~�|����:�or��z�dy�c'���H_Z_n�<��R���� ��I��n�WS��9t5�koY�T��l��[���e����ךB��c�YS�/ h��q�e�y^H��+b�͜�#m)��M�C$.@��^+�#}���/[/k����AO���@�ae���� �ǉ�6��π�.hRÅ�m�x�?�m�

��K�r3�(������>�'uBaή�޶Q���yW��"L���t^	xM�A�;��[�,k:N���&@��L�C*���b�:>�*�2J}~���W���ŋ�%���;�\�L�`?�
��%</��q��.�6U��YDȇ�F�l<�������l�͏��{��PdH|��j4S4Vw	���wؔ��7��ؽ'H򮰏��Uf��<�o�'8U�ɀv�Fu�-�fU�-��Z�~����ۻt���́b$t��&1��C�� �F&�����jP\��R/ ��7?]v�J�}��̀�&�H�<�f��߶$v��׹2�{i�ia[e��-D=�=�'؋7�WG��J��]_A���@��T����i᪆��f�H^'��ʧ��FqE��fffo���Ө�o
`dP���NL���S3m6�b�˜��m&������ih}��rb_�hU�D�fT-mv�'�-0ǘ8t]��}%p�,v9�C�y�fW-����+gт�f~ַ*.�X*��n�Ѣ�0,?J��{���/%��O}?8���Q���!)�CL(=-�ٛ�,nZA�܆Uz�n ��r�z��*�] �!uI[�x,� �7 ;��UΨ5�*�t��#�+�-���թ�'��,-�H��Qׇ�77������BR�:��Y�N�!���{����ܟ�t�k���M����U36ΒJQK%C4��\�)@Q�8�B	�-��-R��y���ڃ,�_Y"�t{\�i�֟�S�ޠOVz����w��-'�x�6R�JL+�A��vj>�����{ލ��y�(v��dD��Le�I�)��Y���i�ma�"��Bť�y�\Ua�D1�2��U9��'2�5L(=��U5.Aq�j>���^K�������Y�H�
ف��{j@b/�����ɐ)�e�d�y�]�G$���6�U��-qG����}J��هvA�>�(,�}�Z�d��jB�IT��������#4�Q�Q/^�N4�1\�6M�/��[����P�`-�nYݑ?��6 �Hi�r��P$�����9�N�#�mo����bi�ۮ��0�H|���"��K�\~�+���{#�C��ABЮ����ߞ�}��Xl�Tti쏥K��auZo5I���%i����̈�� ���w�.k>��3i/�(M��7h��3�����3�� +�dh�Y}�54"���l�����(�"�_����q��b��e�;s6]c1?إ8��)X��zQb��$��|)�_�]�\4
?�?�M9�zL�Mó��Ě��;8vLSss��^"�r�P0f F��o�DS�t�̡���d�b�@�G�;��_��ϡ� ށR�?����q*^/��-�&:��o�ځ�S^Hcz�G��s:��s�]]Q4SV��IN.�h�1�{�NyύF��!#���8�0L�d7�tM��9�!�j3K�VnqI����|]'�A���[�&��c�@�� ���lT��FM1��h����w���T��hM��'$ ��V!FZ�p�.�У^\�([���2h�1$�Go;T�Sp�DT�O�y��b�Y$�wU���]S����Ed7�@������g,=�$e��R2�/��+T�9��!�����������u��sًS8u=�P�X���K�8��Btl��҈v�x�T g�;>zQ;G;�#�ڈp�ꋉ��')�kN�U�MV���*X�s�M��_��z�p(B<EA�� ~�gQ��]����A����&]�؟��#�㟙�(�̞k�ѝ�12v"n\%��'�kE��V_���H�{Di���9��jG��;�W�g�vI�7l�]�HϚ���M��:�) ��%h&���X��
 X��$s���x�}��x��흤:�eԵ�T���c���ީ��`�`�;�#���n��B��7����ړ�(����M+�L��c�aS�sq"���zoK�b�8ygM�Q��U�u(̴��B/0�
�<�I\H�~]�U�1�sSɃk}ώ���`� `�Vz@3�[N}���/#���ʴt�H���`E���F���Nhߥb��2n��C��W�Ź���3�����ۛ&N��)���I�R}�j��XV�����Ya��a�m���c�^����P����cMs*�C����h�Ī�f�.D�_��\ݾEd���L�MiԞ�/���1E_���BS���5����n��O_B�r���Hz4����|�Y�	�'_"��N�v�b����Լu%�1_B���7��iB�>+��9����I��߃��Icd�0����Kd�y6�M�6H�I��Q)�//�t��E �d|j�v�]��q��cu>eAU�G�;7�g6����Z�� ��ޙT2e^K��$���ql,u�����M?4���W��x_�Q+P�7I̅z㤊��'t׍�_��l��갴0JZE�5'��֣��?"�x�>x�8�=GbwR��9�V�)-�>�����WE6�#�f����h?���+i�f0i��fQ��-��N�!X��Bfr�w�u�+����MǸ�Yt?_8�Oi�Qdl:�pSo�L�*u`�=�g��{� �~�����vC���ci���F�p܋��;׵�&�W���5Q��U��1
���n8��0P:�k�9 ܱ/!Mĺ��.�O��"'b���?z�����
���3��7���s���Z�#=�)���ھ��AzD�3s�=�Lgu��i.#3�a����S�v�	��e`���j��>Q/����]��q�9�'�\lLT�+I}7�!�<����ߤ"iˉٓ6�~�c�p�X�1�z�� �~����T�*j��|��ǭ��?�)(yi���"�����cmy<5��A�Z���h���v���c7>6Ǿ5w�?ͪ�k���l9{������W �
��V��� "��g��n�mz�Ď�3V%GA�b�'��+��q$��Z$8����Z��`��ɕ'B�?��\!�}�sq�xx���1�\���d\��w/��eջ�6�1X0�l<�\FLv!���R���u�@�ɱr��`ǭm;ǩ�nk���P�A���Y��9�E3�,��˟O ��y�>h?�DL���yڐ�x��'#(wK���&F!�ᭌ�Ҭ]����4y�Uq��ӫ;�-�m�C)��cǻ@�F�9~{�
�T�7�gC*>� �������F�M}�F.��W]��t;yQ_�巔�� �E��퐟<��'�vwM�x�G�{~�'�p�^ʃ�/��^\]�	�h�Fg�:hvJ����5�8��k��f ���:��H�����k�|�w��zď���5dd@�:@v��	�5�`�q��l����Y��X�������a��M��@	��NIN���7(���F�\���GEb`�%��T#'m�f� Q<w���׬��ԿB���w� 
MP�F��hF�sX�jq�"�/��h�����D�f�Nt�3'k	@�7	�@����*��b��d5���}�����h�g{��" ��,L��`J#���g�ut8Än@Y����|�tx[	 I��x8 �cTdI�!�&�/v[$��Еp�8*2���IpA:g��O�]R�>��VT�L9�w��{�N=/��=�h礅���9��F�n�K�ոe�D[C2�)�9��?��i�������Y?�5'4R�=U��6��=�������Ic2dY���Q�h�Մ2d��0��^B��s�}��taj�d��j�:x^^�� �4]�M�d��'�3�����`���/9n��?�߹�T>�磨�� ��3�'���wР����3���&�D�
w*Q�-������.ZqW	h�+�?��ަzV-_E"ː7���,�2��	L^O��(ž\4��х�xٴ5�O�{k��t��q��T��u$i�ڹX#6�M�;"�?��x'���)	��/u$<�E��brVVH�٪
���:4�Oo&B4��w�1Xt�y<��m��Y��"��Q.�hH)�,��	�\��7�6�@�����؅�ǋ�w�z�^�ɍ�"�j�/���k� ��_$5GW*�%�P'�^�>��Z팮���#xH�?������T�/����[T�\�)��;�noCo�uY�t�>!������u�Q���^M�'Y��g��u��h��=l0ECw�-�#G$Cync��Sǃ�>8���<���Ru9��N}�|�	�v@E���L�?�Kl�%�9��s�/�B���_O�)��J�^�(0����$����[��I��|�wzn�fʆlu��ݟ�
��=x5Xn��XɡN���
��F�
۹�(��b�W�(/��t�K����P���a��!�Xt�Ze["����3D�aK�P�$�'E���J��Ʒ��_]/5]G{�����֢�$#��l���8v-3HK#��zd5���P�l'���V�Ў��]Z�b���V�>�p�L{]�G�P +���
�$�����a1��O�I L1��;��;azn��C��r	a��?AX�vs�����c�K����D�jַͩQ����~$�X���G�N"��sw�F=y��i�>�u�e�X�\T�Q�T�
m�۔�SHR�{5���b�fj�q����'�&j)�;��XŴL��1�����/�lb]�-�<�޼���q@q�r�2E"N�!��T�d0�1���g�._�G�	�7�� !��ˢ�-��;u�΅I�y�*���BH�K����G�<��yxt�p�I�8�H�|�����GK��!^��Qr��	7N��K4A���Tz򔵠�Ĩ���u�D#5=W�hԲ|�2�,��bs����Fh��'�.� r8i���:����3S���,�kBCo���f/�'�H6���`t%!Cb�G;�wr�Y/̮��q.Q���Bv��Wya�hhS���6�!u&o3V�C�����D^x�%W���*Vg�8����%��m~���ș	 ލh+��϶���t^�;�*Lir8��/�ݩ=�2�cQa�5��/8�)�q�/Cz�3$�� �'��L#)%��✎'�Q�l픍���DBP&{¼$�49��\��I������C�N��QN�U��Qqr2v��������Nb�z��<";Jq�T>�s���'͕u��p�{>�DG8,�	�W��z�fXSQa؜W�^�3�P���^Ӆ���K���nҮ~��r��Ji��T`J�7f��k�-�b�H�u�R����(� ����me�~Z ߪ��B`�Ǌx)�C�N{h�mȮ����ܹJ�T�\� ��yt�c����B���pй��sJ")��v�-����}"ɒ䠓�6���z���=M��!&�1�ýZD��1��B�`ĸ�J����h���tt��෱�-_Ö��:�_�/�hP��Q��<�"=�����!"/K�0)F^3Ġ\��#��	#�/�('�ic!�7�����\�� xش�"�$������kv���@�I�$|u��i>Z��RJ��\����ذ��L|�&��H�0�J�� �-�ɬ�]������P �]JiYKc��LV`����Hƕ����"?���j�\��w����0uml�-,��9��x����m*�cHx���6��g�O�#�[*m���q7ܭ�^�h5rE�e�C զ���(r�'��ʑ/[�7�ȿ���Hp}@��%�z�x�UO�:ǐ#�j�1�$t���bD��xxil�n�C��NH���ĠM�����!A����#mî�@iN�s��ȃ��h�2Bk �(M�b�D�a ��o*?��>�1a8d�$@�*�+�'4��r	 �a!p��f���=F@V��5ۦ�&k��(0�Nt�����Nqh�m�1�Ԃh^ٙf�`��逎��5�a@"~�d����9�^�贋l���"e�|���4�@+f����!����m���"���fC���cy��5&/O�BqVٲ;�T5�:�όކ$=��C�k�bx��i!�����ؕ p�kv���D��^�p�_OW��`p9+Oh�q�;�Eos$��W�MI�����K���}��0�S{͎�I�M�Н�7�;˰<��Fq��F��mYg/��)2Ã�is��JW��X+-e1�o�O�m�;�z�^i��'�0�U���6��Ud_�G�j�e��H,r�g��t�ۿ�ݔESp��~%�Z�T�4M���7�h����*���Fy]��9�x��QcOAl�?��l�L��ҭ��ҙ�{j<�T�
�tp:ʕm�9�n%�J-�@�D�#��nr+jv.S�A0/�#/�<5uӑ%�J�p����l��ᩯ���ܵ�G��ӂ����	5N��8�VL��%���#�/>���8<:]��~ �N����]
d!���T���&�(
Nx�=�d�u4������~1��\�S�6c=����㍄�k48���V2t[�Zf���m����%W|���[PE�sIċ�`��KS��6
&N���^�`~.��ґo���!:B�r2fB���X4�_{�+o�%$�w��/�RE�v��#�a���CUc����K��k���5k���!}�Ӹ���$�T��Es@�K[�ؠ*<>�����%��D�P�5�W?��a%��b؜�����2�q�ݦ�;���3 �'���5-%I|��k���*����䥜F�f9,7�..-�Q��D�^�5╴�~طԇS�Jͯ�zl�������]��̙����L���j�=�*�[�O�L��b2ȸ_Dy#߿��Vik�c9I$�!C{%P�[����"o|�F�^�l�AA���n0@&�5����G(�үA1L����1!126�'!*B	��٠B' ���l�C�?� %�5�G��w7�\_�;y�1^,�8��O.�W��Z8#<�ŌL6&� ���r�L�@>hܨY�3O�Ϛg��u��!��a"����ۯ��;��e&$F����nVqD�C�(ϭ�A���wϱE���L}\���~��H����X�qTǚ�fy�%�
�~�����n��_��f
�w��ǁ"�X>bhSA�f�:����w�G�#�)P� �]�$ԩ���wvDP�B/7v��ț�K\Sd���v�,!��>����.���؍�)d�W���A�-p���<}��8IW�.�-sA���o�	�L�6q�3�Ҭ�VJ�9����hML2�rV?���2����(�p�'-��?l)G�%TB�Hك�pFr���Ũw�ܚ�(������2�d�iީ�w�>�9��Q��ۭ�HlaV�E�����	�w����R BA�@� i�s��U`��!������`7�[��� ԓC$��	AY���ӕ�1>����FǪ�Syskf��n��qj?Cq2����B�Z(+2���e�6�Ƃb�d��� ����0����G��ri����o�op|�?�4�ٜ� c�F�X���A�p��l��Np�������J܍�B���g�ȎSޒ? �-� �����wx�����-�-Z�?�Y -������e��ą���x30#���.;�x��94N�㵶U��.��3I3��d9�E���{@�Xsݙ�|k��/q�(��E���r#ܼ��[�}��_=��:���[FF�M�4�ʹ%�o JNFO�Q=3�$8���Y�l�Z&�{^=��ދ@���'���zk�mI�/�*>�*Ҏ༆��!Q&�Ly(ʱF,	���q�PJb��� �˸��[��R�v7q��ְ^i~5MK��Gj�RQԆ�n��~tWm�@U��,} ��F�Jy��FȺ����t�|���&�c��Cꃹ�}�q�ڟϲt ��2����3{�8�O�4�zU�7�@�z՜(��#O�Q
�R�eA3}��gj}�Tܨ]N�:&�k^�Q�dH5���9I����d����'uk�D�}���_�@ed,᦮F���`�ݼTͰu�cnu;����T���W׵��K1��su�4����	I�=�aJ��L~25��n{�T�� �-I��MsA�e;O�2�π�B���6�4��-�m6Kg��.���~
j������}��{���Z�
�g��D|�0R-����Ł�S���R��i�E2��14�B
��<Trc�f�ǰ^�=W*ErRڣa���n$���8�Ƙ�k�����ܕ��r3"Hz��_��^���e�#J�T'f�2� ��NnE^�P��\��
�o��h���'�O�û}�)��M�	�������˘)a��\6u�΁"�>FZ?�K�7n�$m#
H���2����Ā�6/m�I�G۩�<�^��FI�5@�d��2�?��@�vk��>P����K��v�a��?\��/�?�@�C?[+ ���|���2��(�d���[`<��r�/�H����Q��3����O�*�/�{/DeY(��gf��|H�^��aI�p�i?���xSZ��N
5�U���ٸZvf.�?�͚]	������*��^���t0	����5uy�J���h�F�Q�<�Bo�s`�����F�w��t�����1��O �g�K�C�͆����;���Q�1e����d���I�O��@��,�G�^X��EZ�d��+�M�B֍�#m ��-y��eP�W��2j����ʹ=*��6�./=t��u�N_|��dP1����`�I����ai�f��0���9N4IjӦ^�jG��|�~�;-j�i�D?o~�L]#
S��Q�0r�rL[�C��D�?>:����|�Q���tw���\p�~�y���Ҷ h{|M������Nq�{b��h����j}z�R��d��^�nQE��4�~(�0}���0BCX�|eHyvQe�S1Z��B�4��ZOI�[I��f��@@1�E��d�5)	f������[�4j���=7�M9�����-�����N�[�уPL��T�D�_%�sBG~�_b�bA�'� �����4{sI��q�%K7�E5�ڄd�q�$|�!"X	s�2>��Tc3���"9�@2
$��u�a�P�T���#�T�~����t��*�V��a{ ρܰ�O��'%�Ns���/�Р��86����q0c�A��=�+�y夈��v�N�o������)P�9:������K-=ͩ��W	&#��g��*��V��'��N��0T6	ҋ,
���i^�|�k&�6��4�D+��fC�~Xθ�]��y��#�X��l���?��f���뫚}eN>ZK)��)��j%�0�c�1јev5$�Utp��68�Ӊ OP#g
C��I�y�d?/!>�o|����H��:��x��,�� �2�y�F�lNOs��ک/*g$/`ح.[{���p��5;ɷ#��;Na��[�`0n�KdެȤϘ��̍%h.�f��(�ݨ�s"�X �~� ���O3��/�������C�<Ӫ_@f��?/7X���PLMh�nc���JvZ ���:Ѫ'�'�!p���#I����٘��̖�Bd�db�����'���j�R�4$C6O�B�A6���_���96m���qѰ��U�br˪P�2.~c��x�$����Wt���þ�#��3���t1h��մW�Y��4�L��;kBf�վ"�h6��!��Ӝ��,���{�ڸ���rG����ujc�"�	U��i�?7Ǚ�;�G8��f�
悍W}�m"ܲ.��;I�O��¶	�-ױ�⥈��m\>��d��+�Y�	v(S��.>m���?�+���솑K��c������x�F�-��l�	�լl�n?�~�H�H��� �.�!�
<�g������Nd�^�{��&oN*��������m-��\��!P�������#�)7���b,,�lj�0l5�>o-�"�C5&oq4C
��y�%5��p/_�<sk��mF�#7������\�M}MZhh�i�SK�ZUk�&#e��*�3������"
�g���J.�c�+ �j#��?���	���廃!K�"j)�`D�Rv��6�Q&hqc�+E����xJ_�L?�#��*2ǲ,J��S;ʶ��흌�:�����h���-�:��P���QJj�K����v/��?7��Ǭ�2���E* JבU�5��w-^�~;foֈ��cV��ߟyQ�ǃ��������H1H�xJ��oI�U+���#���&�\�a���20�J�8V5M�D�[An��V�`7|����D��CG�Mе8Y��UƌP�Nӣ�D��jT��f]�Ȁ�`z_�l�>O�����a�cr]��z=�k��|CF��1,6e԰�~��-�M�cy��T"���8E�����s0���+�� �a�M]A�uX[א�?�s[ۺ ��Ps�m�EJ��c �?2[Q��9���̶F���7�^�x4�3z�X�t��֑\�H*�<$C�}��h�E��~�%=( ֚�Ǩ�B("��?�S����[�h��	�@��߂�T^t'�[�;Tu�(p���a�O�(5Ox}��"������9��߾�( 1�PWW�}l,(Ɇj|�@�h`�'����lE�a/���,.\{�2vF���ԬX��ǹE^��X@�К��Z[��R�dS�.��
���e~���XL�e�]i��:���E
,>G�9ڶ��a!�Kk��HȠm-����Ǳ��)������+2��}j�u*�
KQ8ɴ�#^�<ys2#~^1�����m�C���6S�s$��bz�pTl����M��ʀ(�A�-`��ˣX�U)
c��D�t�;�r�|��g�v�BF����M�Ȳ�iY3�D+���J��$CE�C5�ǎO�g���W\B���Q��ӟ��I�A��D~�tx׳��kc�~ԯ�="�	���e<T���q�^u�"��M?�z�,9rK7"^��1���~�-ŷ^�UtЙ�#%t�o���+�+�0��|(��E����j����#�S/�`�n������3��1W��+�6�"�
L�G�����0�3�|q�wⱿATt���}���٠|��$��]��1��?�@��x�ṡQI\��MgL[�����R���B��7i AN�\���U[����"$�Pu�����l}�JN�0$���}Dx!K�	zKg�v*n�O�'`I� �t��S�� �H��J"Z��ܯ�?��ؠ��:62�.���ܱ�]��ϰ�5R��` u��PR��D�+�G�b+��sW�#BX��G�}NA�<s	b<kr�%���7U]�7a]B+�yR���HA��Kƫ>k�����b̥���c�O���GN;�U��ř������od%�X������R��'�*J�,͖@a&�.��y�\�/��C�� �}1�n5k�wG�\5ٲ&�V��gF�p�S����w��F1�,�M� �墒wKK�5W}�).���ⓢ2��yȪ����7�8-Uj�E�y��+������M5�O�
�0=���&��o���:[�=�q�ӑ�=.'��g�M�+�2�/Z얽F��=�|y���*�ί���R ����1jb�BZݬ�Z;N
�\?���X�f�S��߭شWԂ�Ax�fh��e�|7�HX�最E�w�qY�,�7I���"���r�o�ܬ�;�]Y�������HkO�];GT��E���Y��(Ή����%����+�z)�-���/�b�k,��s>&_��gx����tB.=Ni��a�f� (��
�F�S2���;>ۓ��r�y��}���D�p$S��Ʋ�������%�K��G�'��6�|�X��C7N��]̣�S��t�����9���ЛS��y��ˠ�}+�,P�b�f��uWE�4),��"��F�������+}�`;2�֓��P�55���w>?N��V��v��(9ig�k�G�z�A�	�~)�~�&[�;_���w�����UއQ���J��	yi�m���>�a��Y5Բ5�65ݤT��x�H��f�@+��ȍ�b��%�,"�QF��W@=2a����*�m���F���&�
ܟ�U1���2�c9���G�"[�(j�j�K���F����s�3!��m^ĸ;>|'����K�>3���o�n%�䬓<���x��!w�qܻ�5'΄�,�H8#��34����f�3Kr�����,�	������{�hOfM���P#��p�)�L�T���G����tB���P�[�W5:�@_��RR��5pw����G�F�qJ�5g�J(� ߭�nu*���^���hH�:4Y�Ԟ����6�:��YzӸe��t�+^�iW���̉���#�S�y��-sg_�J�� p���e��^u��wH�D�6Ms�A��-p�)CA�^y���v|�;�<���!���?��������%zu����t��^�����ߩp\\fJ�C��@�E��x���l	�+ĭrE��e���j%7��|_7�_�N�_w���8F9�\�p�� ������`�]�R��A�Q����b���ᘀ	���R�}y/�p�>��Bǽ�#V�w�I�IK�\L�-���Z�*s�d��zy�������{:nn���@��FoH�q�-�F'����k�uy~"�(m,E7H�.��z�o�E<���ɭ���14�alAQ��@ ��ы����j�U1�N��^$�'�m��[53�4 ^�~,���F �dC8M��c����ˣ���aM"�j%�I~��X�y��\Nj��>c�@f�L��=p2�����eHw:0:�t�}�,Z'�IA��<�Y�"�(����Y�}E��E��W�V�1c�V&X��SaˡѠ�g����5������$�^�t���F2���t�<����$T@`&�8�^�.2Q�]J��N3�ZQC�������տ�,{C��ǀ��H#@���9�\Ø���s.�����Pp���O
#6��jݹ��孨!��,�Wv2)iY�n��=�I�iP����/���ү�6�LΖ�����b>5yE{�RO!D`5��g�i�;�X�p�]�]ˎo�P�sfNw�A�����~���U�5R��g��."T}_�����:�kq=����o�c�\ۮ7Q\�%6�Һ��+)�F;�v?S�B(Ԑ1�7{i�c)�9-�&��w��g�L07 	E ���3:N���Md�)~��
	�z�-�>���5P�P��9�Vь>W��{�?��-y�I�[��E��~��-��C�Λx�p�gͧ����Α
��f�,��w�E\�H�~�b$Lp�dB�{�.�&@ӗ��v���n@�1�rzo����C�ԝ?/��6#�ǔ�:��a�@,�$-v�ʭ{	����D�Z���\�h�O���$oO���hn%�dVxP4l3�N衶����J������a���rvc�d()�͞^�X���r/`Y�nG���,C��=�
J��0!Q�?�K�u�����V��C�(T����ں�X�S�9d�d�
,�>��Å���ή|����s.I��P�~�p4��%,5��nNzm������:$+��ߺ{��q��o�k(uSni�B7[8@w�p���d��W!@��k���u4[b��=�D�|m�߹jmV��Ր!�8�#�vhy#�X��X��*��ʍ����0�+�.}��9�v�ʋz�%�棆��s�Q�ǒE�XiņT����j�9"���e���_i�P�k����N�oS��"ć���'&^
�A�}���|u :�>99]���M?Ԏ���O�	�y���[	�D ��C>Z�ӎ�+�|W���|@С���4��j?y����z V�	�9�`a j�������b�/���6��rFʴF��MMU���6v�Qh;�p'�MEя-͸�蜚���8�ɩIk�q	0���0� 
b��պ�ɏ��Ō�~��xwk�i������}bg�r4)p�ʓ���Ry��R���,�	疎ÑK�Kݿ蹨���}�����ƨ���U��-}�N@�C�6�3[���v�7�~c6��P��ӳ%�m��`??H�t���
S�5�x� A������?,"��j���Ҭ�-|b)�a}{#$౿��0���p���U�Q�%�2�����<�PӃ̣?�1u�Bt���,h�5�:�۶�R|�j�-�2:⑎��V����%R\�6m Վ8�0�P`�b����c���Ӹ�DD�����*&���/k�E��X�i��3��z��@�͎Țgg���ܑ^@?/u�<�7��{c�p�S���bo)�� ���ӎ�r^"�hf2��������Gv*s�Bdl�c�� �r�9`���42)�D�ݾ���^���B���n3��W#HG{���ENe�v���\��j<�3�.;i�>���i��Յ	���&��j��VQv�yG���q���r��τCd[Fa2�=�6�ւ��K�JSm�K��)�]Α`�'r�;�=fCՐ�G�%�;?�`A�t�>��	���ӹ�YWV:�>����|�!�_�Q�ɐ}��I0ء�d�KΨ���.A�j�#~�>/8סؘu�gX��u/v����>��_tR7���+���"{�<��z�N��F����z4k�����ST��9�V#�H��ZK�S���J��|�F�Kw�MA5d*i�Vc	�%_/��>�4zg�z��2�:��}G�����ϡ7!�PP�~A'4��Db��!y!q,9��ԝ�~���*S����ym��a,���L�l%dV�b�Z:������D�����S~�E����e6ʋw�C&�a!������|jj���,���G�U�[;}���	�h���?���R)t��V[�F�{��R�/"�H-��%����k�J��G{ ��SfGù�F����	��>��keC�7��*f��]��{qWG�ړ�a�V��3��	*T��n�Ch� �|�3����/��P��{y��hA��L���Ed�5����+��2����c����������#��9�#�D��/@r���r�;#�ś��u�E�`�[�%�	+3�d�g�-pY�z�х����7��P�`���qM�6D�rg����̮��z^ꐝ����7ц��	�j'��Y�+um�I`Qh2')�ƫ�{~a�Z2����6�jٙ�0�up�a�"�Y�{7��=T���&T(�����ٿS�;AП���n/q�Ayv}���v#�{`�ؐ�H���i+ӣ���uw���u�V��S�i1O5�L_f֗s��kc�D�7�� Tj��x�$M�,(�D()*_Zձ�#1��ބ#@6�'s���=Oms�b"�=��4�:�����a��}&�Ed�!cW>"���?Z5��T��g�����\��-�Q+�ĘkN
�k"�q^��B=�q$]��@}V���wɇ�iEi(��JVa��|h�R���t׎��ǔ��
�e�v'��c��눅��?W��d2�g�5��=�Wv�Q��_x��}���M�4\MG�φ-	��hEC�j�]��W�P���;�@��Oc'ax_ �0T���0ŉZT&����E�#�mT�a׵K��J������(>�f��B���8"pU���}#��'L4�g(��C���=Wӕ�\�v�Z����2�B��� �V�[_r��h�]�HI訠G2n1:�x~�b!qe��s?�\:{��t�Ex��&��vp�$D�����nu���A���+�4^ƼD	5�)��1#$j{�>=�~x���l�K,��ҵSgW�ד�h�H��(Z�(�
���cm����31��%K�}Ƨ�s�k
1���{3�E>�K?�UςZ��A{t[�O�W�����G�:�����{�Z��N_wt@������X+gF�Z�N4�r�R��Kԣ�t�vw��,���Y����U��74��u����(EG"�v����J%�x���¥+ŽI��o��B��2��"As�S�N,���Kp}���U��eJ-8��3�*!�y�Mg�	�F��o*���[���� �d�#
�G
l���FfU�[Ʒ9���_�H�����LH5���P���dJ
�X-o�Q��1NHCuA �a����q�&B�G9�Xd��(�s�
ù%��Rړm7~���+ ��T�G�ɏT���*��2�d��\�2wT�Qt�<�����;������OZ�֕(&a�Ov�#���,32�U;S�t.p��^�x�������Ŗ��$9g�g�Ξ{b����!�H2�̶����FQe�Q%*`'׫S��܋�#��NC�OS�'Jb�V����9~6pAq�^��t�W`(���*ۼ�Y�
d�e�;��h�B��V�^{�X�`�j�Ď���,�{z�럟@��_R�G��lt^�j}z��(~��`T)��B�_�r��������w���9�0 i�gDH�K�h^2�f��	�M>e�Y�o�q�>E����.�>�@�x�p�F,]&]���8IM\6�}ڟ^�/Q���� �Ij*�^�?�!�ow����ϩ'*��)�J')�Z��eџ�S�&��+1�hW�D�����\`��1Z���Vi6*m3�jNB�ʰ$��"K�Đ����j�41Hd�C>[!�^c��W�-�&��!h�:`X0B"]��+�/�D�鍗�)nl#�2�b���6��]l�=�����vǎ���_vLװx�ŕO����Rw2�b�Q<�#L�а����|*��o�L�1�C���^��-q���?�m�[MvR�&��vQ1ab�:ئ񗷃�h(��T�`���H�Ġ6�M��t�-�!4���-r�,��lvh�1>M݈��g1�=;��� �A'~�ayZ0��3q��=;�7W ����9��/������_ ��Z��5�f��P�isA�'�7^:���X�#�'~g����]�ʐ}�;tw��k��:��]��?���
S\���h \�7�������mP;��L�
U�<���&�A�LV֧�Vyw��6ס	���+����w�\x7;��T��,"f��ӹ�_s2���)9Ua����m[!��j'�_�I�d;�^R*&%�2�6EYpzQbֹ]K'�<���DdZ�ٵv lg�RҖ&����a|�"䑸�r�7���|q�ňU�O��i�ll�5_Q���dbX4�XLl�*�`F��,�^>�Y�y
�P���=��8YG�B�5�1<��eQ����2������yY��u��^Rg�LC˿+�l_r �Hƅ"�FN�[�l��*_>�M<�QwD��1�gN�"�^���g``�\N�<R�<]oU�����EM�Q`Q}ٔ�=��슗�7��?Y���=Z ��U�1-	5�敢<�o�yEA�CdƑ�_���υ�QtW�UFO	�a�K�sh��E�g�̈́��t���_�UB%���s�F'ǫl=B�U��ۯP���JkF�Ҽhi|'i!�AWŃ��}�ة�U���Πe^�DP���POѝ�cKMM�Z��TD2Y_�Fn\�'5e��g!���p/������N�e��0��N|o�V��L������.2�޵v���S5)kz�����S�7}��m�H������檴�w&�p��Ł�,�����I!޾Q�g��3���г�{�;;��Ğ��T�H|i�7����k{�\̩�=��^WR�!]1b֞�E|�I��1�Iv���AAvn���W�YWZ�Aɦvj{`�9C��5_�E�I�m�20(b2����H��{��ͺ�J���v'��y�d��������ĵyX��A�JO��O9�2���S��M$�p��Ҡu�G�w���%`���*��=�u	# ���Pp{J��se��!�n�%y<r�Z�y��]bK�'N��1j�׵����� �8LE�a1��Y$`����
�����T
�߁�QLy�;[���4i�������&���WI�<&hk�zu�`Lꑲ� �|�a���|�
�3 �91��@��uJ(k�='.@o�y$���J%�c�#]���[��c3-��m����s�zج��97����}�'	�i�R����(W_ ���'َr�S-��S��a�Qp�0��>��)ke�ª�~%�uM��Ź����Τ�\��!�_^���a?;k�nً��V)ϔ\9`f�ʞ�y�KEs��&f�L��?اd��:7<��t��`s�<��x�{
JL�6fd���Ʋ�1�ž� ��"a��!���?~�C�VYs�8zb�k#�G`��B�����zO�z���(�����C�gb^[N�!���v����+���|�$��ɎU��R.I*� ��˯��h$2�
�j�tw�Ű��}TN8��a:�Ģ[E,�W���YC0Ȳ;Ķ�>M�'Z� ē~�$�(Ӗ����6: FS�6#�O��Y����+�^1�c���Q���e��m.g@��95���������Pk�	�d,K���b+���Md��HQ�?O��TOB}��������\�� �$�|�" �6%4���z��j �B�*e���]N v��K�	�2GO��-s��&aDf�Kb�By�ͭJ`�����F�A���i|���^$D�R˙c�jLzH�%��� )"���&��ob�y0��J�;c2��:P�+���E�W�pG?]���9:_HM$>�Q8��-YU��0g�Y#�kc!� $Sד�A'0�w��C4Z~��܈�"0��ٻK��d/@�Q4Ʈe���U�����k��LA�T	\�r�0�4�@���q7�ka�|�4�P���=l��d��;�e���^��.0�t��g�
$j\:H�G�䲨˓��X�
H�[� Z���Nۦ>E�Ы�K�P��ksv ê���H�e�U������LD*'�Z�+ɵU/��~�:U�C�;6�v��-��:s�ڀ���h�;n͌�f���<ٗ��g��\������F(DK��RW�$�-���,��k������T^W܊�<D��ƉH2��QkP�9,gz���g�5Ha��$6�W��S4A[����)H��< �����do�H��(�{����u�:Z(��.�g�[	E�K���0u	���2��SiS$oU��487I�{�i�@b�Q��/�n���e2`=g6���i�߻�r�͂d�L�C�N������M���6	1�/����ū��l}���"�B*˞�꒏�Q�`�-G�<�h�?E�()�79w�Q��r�mD0C��������oƖfB��Ҙ�X_.ΆH.^���뜕69��/-�GW��n�L��o`
j�����L`�/o\C���[��ԯPD�r�:n��s>pb��?��@t�a�EAf�W�[�wݔ��F�d�i=�V�uh����Z'���VW';hﰭj�\X��(��h{F��\�D�����/E�kJ�FX���ڛi쭲�$��S���S��SI�i�X�D����Ʉ���s���9����g{��b��7��.�04 �I�����M��t(����c8՛^�W�eE��+�B����ڥ\?���m�<ʚ�� �
Z1����|���k'&3�A��T)�?&�q��-�(����W��i�j�����!T�4VH���hm��Bˣ1��