��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c�J\\! B-�B�^F;P�sοұ��z�Dl�~�����u���?T�@��ۓԭ�+�{~���a܆5� �0ChY���;���6�Tʽ.B@�0�B�޽����>�@R�s�6�|Ҥ�
t4���_*���ׯ$�ѵ�d@D���L� 9}�6�4�H�u1`1��K@Ks/[�-���n�����o��'"�i@�m;�۩+���D���agA��y�R�-#Z$j4M1�raX�L����v����W����_��V�m��饵�#:4f}Wqz�~��D��:�ǿ�WUrG^���Q���(ˍ]�&���H�ØO���o��|��N��#)aͱ=��6́
��qƓ���\1�������/��  ��!�F7ݔ���1�J����4�?�@�'EKG�]�40%xDT�Nt.w!Iރ+���Yݯ�����u��`�k���J�S����h"RP��c�u��Ԩ�Q�`�*@ܾ�7K(·d�$*�h�롭<�Q|�i�� �K��-.�
2�x��,�TTP0��3H�a���SZ����h��`e\BH7>
�N��=���Pg�{�0��R��XQ���n��{Y�G��Q�N�����^<�R��^����W��k��q�XbD�~f��6��,���Ր�7�7��$��k#�gm�]{��l�D�	gq��j�c��w��3�R���u�B6bw��J��=���6~��:;�8G��w�OeК��o>	}���wr�NX��L�j�QL����THV�LJ��(��*�U��E?�6ki������ $�?�*B���� i'"������`x~�X���OL��D�6z�V����	2��a��7�k�Ռ��0�1q��YM�-0�Pbz���O$I���Bճd��6�ml���[V�)���R���C����[QjEp��$l�����Z�LNQF��>�[�36��8S��t�pm���$>�X�h�V����5��5���^����}Hϳ�<XY��<8(�f����C��鵉t|)��P�[���'�w���"�����:V||����Y��ԯ�j�)���i0,���zC��A�yK�#>*��꽅�o'$ZQ_�'�<W�w����"���_�ܸ��7CdTFȁ�$���B�q�P��}ո~9`��얤��`[ӄ	���n
��/pp���'�Zh�z�eQg����|�*��5�frB���]������UȤ]�I?1����4X��w��n�̳�Ĺ��/������Q�s�?����ȣМ���꼁#��&��JO�� ��M�̻��@i.�� I���l(��Y$J$K�J���#�Q��� 6#!��G`!V���d�~��բ!lC�����+B���S�g�0�ϰ`]y�&�
@�t�cf����t��z'<��`q@� ����=�LG��S����.���S��+�:L�_�Y]w^���ԠG9���W�#.7oB��N��ҿd_Ǵ�I⨻�P�.�j�Օ�E#�*��K�,Q��7����ӿB���$��Hb���o�ҟ����v�S�O?.�[Fr�1��b��o�="A�d�@�j���j���`ӹ��)G4xq�2|��c�ƶV�6�(��P|)p�7�h%;8��21���t��(��h"��vpO4<��Z�q��
lňGѲ�hk%�0qu���JS.UYb	,� ���\�U��h@�v�柢vUf5���L��W������&V�V���K��2��V"�7�  ����MbC��z>����Ej��+�
���h^R��U���Pv�L$��e5����o�J�����%>�@���QЅK��3�/ ���H���}�|ǉ[�q�n<~�J�j�K���F���E5��J�p��y~ز��A�.I���KU�W,�V�X��x8VP;��q�ۯtJ�"~��=����1�|F��;�)�K�ǐ�@���f\w���5ٰ�Fj�̠h!vPUt���¸Գ�,������^��܇JovB���t3�����Y��x���u�p�;�;c��N�]��L%:}�����ױw�m:�"��l�S���w|B���q�>Q&.�5Eu}v7�;��lb�����;���X��i��ͣ�U)�W�Q��o�U+jk\E�J;��N�E�rs㥍�G2b@N�1L���{�QO�+��2 ����!QR��T�*����$hr�~��� )���s�k��{�ݓ<#�:f`�R{�%HC1��?�S��7;+�`C�^3]����(��6�����g���k+�t�D��`��%q�/{~�a�b�.�M*�?�<Ri�e)�-���$BF�k�c�|V��.^̷�Θ�k������$|g��f
f >I+jFU���GD�:Z�l>�*wg<%��*J�������y�Q�~)������Y ��n1����.Hk�㜜�S֔ߟ���ˑ���*�	\,�����cv�J�K#?�-��u~.X��u��I2g՝�[q3A��FegU��a�x�S�f�AG�A�'�f�*8�q��
�gz��$ɞ~(QpG|5�����E���� [^��^ٸg���+nM�.�I�4
k�u�D!�/��/M�!�U�Vʟ4�G`3�ڥ��zC�J���^�&�dh{p�����Xy�0&ߜq��V��}�Ȯ�$�ZR�L�����4߶������P)s��"l���6![�� z�[Ѷ�/��%Y�e_��n�!�y#��2�3Wd�R�� .�K2pSߛ^Q^�3�bS�����#�����˃Q��݃n9.��]C;��(ҡ�Q'��V�g��۱�f�[�L]5���&΄��|1a���֫���GR���Cy�+�s�:[D��k�!(Lq]��Q��Nw�E���h��\�#�y�B9�Y^�cY�U���W��7pF�����;6 �{r�ZI�ϱJ����c#_z��K��I�a�pH.W��r�W�'�ic@X!`������t�[�UyQ��@د˓�{�?{k;���s;"|����< ��E������ޥ�|�S����=�0�0���^{T�T�����,�����R����b�2��;W갡]̍�R���.Ӻ�t�*������ҕ��e_��(P�6t�>�V�5O�S{Z����w+�VPG�&9V+W��*�(�Uk�d0t�βH�MrM�Ky��ɏO�V	��'�^�wv��o����+9�Zc8�Efo��v!���²Wȩ�+���mI�����ӰV��F�[%����u���,��-�׍��R�?�s��1�+�	��hLԶ]��d���̴Po�D�{qjAu��E�Rb4	�W�OC7�2o�P�v�w�!�E���$h������B��f3d�K�5��6\uY0g�!� ��}�������W�X�L��O�"ԗb$��ll�˷'0Ʒ�<4v��y�X5�"Hɲ����(�^)r5�A��G�8v�J�hR�*�HQ6�̦�v���	0?��9�<ݨ0K0!�����'���d���&�<�\C]L�������u�6�~�ҐI�����B���a"���TR^E +T=/��[��7h��0q�(ͦ�L��%�=�I�Xf.�g)��i�]4禗�R<hoT��K��.;�.��3��C��!�|��6���-��0.i���,�JԬ�{���^���!�V;�o�D)LVv�t��tJ,,i�2��ըS�H�\���>e�C��9�+�[מ�ŕu�!L�����n�Tv��@K�/|�KR�fz }�
~�|�AQa���i��P�H�'1=�\��\qi���6!�)�d�a�0x�ȆÙY�b��5J��G{d����x�wt0�Ab�\�g�Vvz�CH~g=�
aYFa*��L�y���񍣳O�/	Z���v1e�1~L-�z��PC_��;	Sd2�N��_pz�Ŋ�-���#��@��%ʓ�	<N֙�*&�V`E����e�"��T�7@���[�Ou�!�!�_=�[��-�^��,U��ì+���.�~IsY2֧��&�Tt=ޡ���jf+O�5k��5���cAMؔ��;(o:��1T�
�u1ޘ�D��V�ո����)�!A���3g�#=�%#^fs^�s"��H��#q}�R��UR����t��I�YMBt���CE� ����K,cvD�%XKj:�����.9�#�~K����jS섥mN�	35 `z���3fc�I&n��h�L��O�+~�mj@ꌥ�8������ݝ!�L=5���䥠~+ثq�.O��?u�e��ǲ*�X�����cg�0	S�dbD��os6�K���\�(��-�{iJ8�6���?ޗ�u��4�R{IJ��Yk�dkk�6ıH�+�;h5����9�M��,�!���8(.�x����%�^Rz [�Y�F��@8��N��X���ʠ��-z<��-z_�����̻���i0�cP�ei΢�r=��ep�A �H(6�cDvy{�����D�$	'���wR��J��y���A�;����g��kd�[�6�Q��X-�$ =�	E��|x�kn���B��V7N^�]t/��?��j�N�GK��,�qȲ��!�J���WYXf��;��lW͎`�G�1�{$[�3� ��"[5^8�%�� 2��D�!$�t;�m�j�_�+��j��E�,��>L�#ͳh��k㍯FP"p�,7⯱*BT�=?��4�����(�2���;��S;#j��G	�x��HT)�tB�����/[b�ČY8"wifY6ߑ��GVۼ:ɖ:l�~Bķ��t���԰\�K�����b���t��̳m-]˺p��>�^�����n��=�/H"-���[�3�x�:j�����4*/��K���<�(Yrx�g<��y�Í� u>��c��P�}�i�5�N��-z;	S]im����P?���,�^��Hi� ��:n���5�-��n�����Wr3Ǳ����[1CG0�?��y� ��n
*��u���4�%;����Dᢖ�Qg��E[�UA�i������������B���<��~ץ���#���=>Oy�[	V3���ʿ�A��5e��#���>����R��Q��t��
���'�\)φ�DQ�MD���78�r���l]������bӋV����O�����Y2�6�>N^F�d��$�Û56����DsD�N���<���E���"b�W;w��!N��Xp��SI~o�L:G�A��O���d7&�JՅԶ�$ZHgHL��z��u!�rP�)m�܃�k_�أq7��ƜN�Tzٹ���@#������J�v���)�T��M�����~�?�7�*x{���jћZҊ������g�{+����J� ��$=�0Q8��gF`�?ie�l���-V�LiK�Qa=Bʎ������0��\"%_Eg8	��Ӎh�6����A�z(�KG�j�4��N_���c�9>����VǛ���[�C8�Fq�,5V}��w�`�� *_�.ٟ=����\`H�Ì�z�+�j����5��W�~���8��׿��:�JL�U����Y��ʙ8�K�?�b����ح�Y��F��h�z_H�6�ƹ�#��]�</�͠��5]�q��u�����-ލۙ3�6r�/�ɡ�\����c��ʲB��{io�d��%\����X�s#�^���:�4�[���B���L:��w��?�Y�
(bkk�=��I/��1ի&���E����"n�7�����Q�ӲWϩ��Y�>"�j��桯";��#�W0
���x�7�8�m	K%��e-X�My��]CY�.*�ŀO�h#���X>o>��щ��ņk�G��ll�ºM�2�������	K�4Fss�(�-�A"g���c�_��1C�c1��+�Ш���_�7><��x��j!�/m���=�#ݩ2'ә:Aq����ie�YY��Igʧ����Gy�3��R�]�7.���G����:1���*Ī���h�����}.����P�$7�MB�ٖ��p�cҔM�ۂ���NGaŒ݂�Ii���a_B�V	3
$y��o>��t�X93q+����������N+��`G���@D��hb�"~�9��ȅ���V�%��O]h�ٶF� S'�q'�S?�p�/!W�w���U8���b����j���ktYr�B��h��YaQ�Yl�I^��	h a|蒋�����j��w@4�]m�)Ѐ���AQv�����%�y�r�R���L)��	�y��TZx��@��(ulf���-TU�Y-'��e~?�����eZ�~��������1�����J�q.d��ew�2���!��n�MƸ�B��eH�0�>��Z���5��u�AwaG�O����(�����*$�� �U���'�!�5|����1TTڅ�p�<�Aɏ�S��X�ޚ�_��/��X(���6�d��eUmj�Wr4��Tv@��iOxh�����rݖ������?��]���I����Ċ6��K���[�aw�)k���d$OQ��'֥��U��/����j4��qM%k$��M��h�Ql�=��t��>�Rj��^[c�T{��_�k��s�E�掻�)�^�A�<�}�h�6�������e	i��\&�@}B����9�XΗ3�&�۵ ������J�d��h���)�X���}�X?@u���6����h����[���_������� �+�c�]%����/�'Iq0�e�RUbD'm6*R��]�+������k'7?S��B'_��к0�� aπ���'oh_H�>Z��&�˯��>Q'ݩ�#N����;C��3��:��a|�g��:�Cn2�>�)v��zO��@�&a	V	ݵ��v%��B���p8#<�L3��jN�J���D�}U���tQ�Z��
��w!��̴�k����vf�%�#�F��/_��rվ=�<���������"aHt�1�����1�B�f�yx��`6��*�(gF��o>��?��0lF�D�(NOPNZ�:��σ�6{$�:��W��;p���G�}��d=����iG}�y�8����HyHLΖ���_U��.X�#s��Y�����T�����^����i���?��5�N��H�u=��&t}�n*��vӸ�L���<m���)�-G��_B{��A2pw��%�%F���d֭�W1���S>�6Tb�31�OOK\��Io��'?�ǀ���#�~�+�{Y�9W������o��z*���:����*��f�X�^п3�L�tc	1�9���}x�L�������w�spc�Q�\�]>o ! _C�䩀�CȯXS��+_�ϒ���9L(>)���~���}��4�]�Tk�e:s
���/`
(�����@N5�s�R6�Ld�Mq�ƐIKr�7)Њ�õ�|���f�Wjko�&�J�uc63��hʔ�!�l���U��ݔ���ח�V�ͽm=l�6�~.e�1�1ɪW�y�]F/vj	�/g�S_�K=�S�)�X	V�1���=��r��L�_X}��l ��T�
݃�&�w0�r��^���i�C]©M�V�B�71�9�N���,���WC?&O/G���΍�[{�ֵ���3l7[�W��y�0���ԗL'|��C��a�Q2��u@�.�3F���s�r���\�����@�����'1Y�2�m&�i�(*������f�L���DZ�,���J�o!���N@��㉢����;)-	H��D�˲�cl˔�OSk`��� �!�쮔��{�2�P拞`��\5	��O ��t}��������eQi��W/ev�+u����jʽ��W����~�\rVs
����FLv�m��q�����C^�G9j�W.��;4*��9(��p;d�<V
�P���]v�QD��"��Zj����(�X	=K���$�_��|u�I[�͌���CS�-M"���p��"�W}�A�Fp�rɯ<�v詍:l��`���k!��*Z��������s�'\n@�����'��d�@���8��f|��kœ0.W<R-�K4W٥d}�>��Ժ#B�"��}C�)_�e�6_��"��J{�����L�2�����&Vݛq��ۿ~`;Q�rT�Z�q�D�c)����7~t�.�Ȝ�?�7�?�� �-Y�f�Hz�"nح�*�� m�"��̔�r��-p N!ó>L�ut�w��������U&I^�g:�V.��)��L"��=��[ N3����x6&��	�}��Sx"���p��Cnqi�����{#�R����Z9��9M�ַ����x#.�څ)!GV�Wd���V$f*L0vJ��S�����t`���j���5���s�kl�lgh[;up�L
G�������0�5�檲3�s�u�`�2��^�}��Ɔ�;�D���ғ۬/Pe�j���`��.q��O�`��ձ�$���w�3O�-��z6�U��=Mf���<H�{�a�<��B�M̿L�\岮���@I��E�\=��½���<��Ҿ�#�a2���\�?�_���T�g~��r~
��al��-�����6��Q���@��ٴH��=g�͠�sv��V/%6�����#�Q���=�&��a�ƹ���}]s6|�1l�<)6�x�U:��:�܄Tb�H��"�/�rQ�=�٫
�BE4����RE��x�y���ρ҉�G��[s�x�ՔI�={M��E;H������{��[ϴ�}�n�%���؉�F�r�Ċ^�GD	E�����C��"�w�I�o��E�CI��S�V��}�}�9\we)��hC 
�KC( �Յ�j+����>]ѠDRӡX�ھ2)`�w���(
+�Nh$S?V*��u*ܷ�T�`���@�OM�z9��r�V�J	�^..*m��el�p�v�Ҙ<�S׽� ���l^����} ���ir�� "s�'���3�CڎW��[��DI��SxE�ܐ�c20��|���gL��(����6�h�����P�J�;�'��eѣ:��L�^�vU_�j�ʹ4��r�T�6,���D�V�����릣������������/�4N�ge�>�_Z�>g�6a��)�F��l���	'^x��A=AG��4:�f�o+���5[�>'D]��J<��08�����Cq�X�.%Cq�J���ξv.^ZQI!/�����z�e��Zzv���&��⬅�%�G'$�źţ�ć�!ֆ���Ί"~M����CT�+�\/<��/d���?Nu<�8�Ұ�8F2�{/+���@�͑l�?C�,�� ��0���ݻA�6 8i�\;Zv4�ڸ�̲,S����~SM }��P�*m�3�h��c춧o��8\\�p�8.ͳ��^=�p��#�Z�C��'�`������+�/U0󯁌>Cȉ@+�e��7$���K �J��T������h�T�����p ��V�x����0�!Ő�H�����S�N���o7ς:M�xI�Qn�8&�V9���%�hF��p�N���y���N�#��Z>�0{>���/%���v��L�I7
!s��j� �^����cտ��6�*ÿ/i�rj��og�C4�4�����I^�Xi.���mTޗ~��>~`�?�Β��N6�܄������TUp��0�5��	M����Y_vF:�	٥��G�{�N+7��!1�/b���*�i��4������l@z��q%$IԲ��"�%1���Y��'pzg�g��Ѳ�.Bb[?�EǊ����q�4t�c;�����,3o?6y�[�V����a�:]Ķ�(@�b����J�݉IT=���R���u^�+ۡ�O�� v�?�Jui�yɍڀD���o�/.� �?���)�'�f����H��vGxY$�rq���@QWև����{����b��@��,~�IK��������J}���0���6�78��x3���]�ƃ���A�M<h�T��;����z;{�߬G|\Iu�E#�Ke+@�<P�� ��]X�e�U�j�$��xj�вOn����!���搽��֠�v>��H��r�7f��a���_��@6$*���-�ŕ�\�q�.�朣��sX�z��\���a���B����-�D��u��~gs$�l�Kg,C2F?�5"F���$Sl�2���n�F��s(��F�	{(F�������h��K��N[28����+��(���-�~<
5���	��幫�h��U�*I��~�TrG2P��#�p%ʤ+�\�Q�D��Ki��8� ��jwv1kF��J<�,Q�U�m �G%�_4�������Q�"\�����r	�Ч�%Uk�I�5k��^Z���9�=�з�E�9�"J�YH�%��L:q��,u_��	j�+�(FČrFA�K!����֏����S*�3�,���o���_x��#9�� ���#���熥�V{�w��n�ܙz��H��(��Q8��ӿr|���{�I������ ĉ�!჻N?��i�ͳϴ����#Q9c�G�wJ�ik&��+��w��W���L�]oq�_�-���0��ܒ�p��� �U�� �����{��!<**g�#M�Ƹ�ӛ�ī����Nͽ:^.�%�A��o
�����D���㕴���k���S�u.1����J�G!�9����Oe��y���yE�`眰\�W�4� haH�U�v����Q�&����Y��� �Hmq�e�ˆ����?�wi�"ޭ�j�/,�0/a5b�(��R��~RȦ�Je����%���Ҝ2SX���#�hj���W̕�Fc��~� �H׿ӎd˥�s�Geu���b^�ն��;���ʼ�n��F�$�o?ޞ�`�g>�����J�Bim����C*���SYa8ʿ&ޞ�taG�j�W2�r��}i�*\���RI��w��ZޚI�\9�FI��.e�k+G�{��]���)�݂��q;g�iqU�xC��7$��K�{m�d�ݠ!�h��d���l�Թֶe�[�"���1��6�ɥY���L%q�n���!&�p�<�/6A��&N�� 2�S8� AW�oz�}L�z�9��	��đ^����6r�f+�+�N�V߸@ �FnAk���.��F%��UxW:Ǟ�;�u����\����g;CrٯI:�=����_���T��k�h�E�����f�����w�+GLd�l��'�Ӛt�@��+1Y��:�w��rE��p#]�9�k�Hnl�_9b�Ml׳��i� � �xʫ�g�*Wօ?�<��֨xrz��1�����o� �=��L��]` w��>D�1!�G�_���	-,A�'+=�$N��75��m\`�m���������\���6�DF��%AƜ��L��҇�X���c�Ya��]��yw��?���c��v�K�7B�ʕ�,
�����,a��e<���H%�Č%�ܹ$EN\*���$�Jݘy,5�2{�<Ϙ��kcq��a���T�p��?�vr�������2q�ѵ@*0?�n�O����ČrA��:L���E��T���b�R*UGVa��I�����
�����i��l�������Q�� �]�@�@V>?�QM� 0I~��i����ت-���ߜy(Ӯ����lew���L	����q�Ȓ6	��g���h�$-�U�3�W�nH��@��L6��n��k�"�7�/ h�ޑ��YTB���CPHu[������ G��=t����kp@�Go|�ݔ��E�1�������Z�C�p�d[i1-��P�����)^f�l�4tv�V��w�	+i��j9�r8���	G���D�a��)V�J,EΒ��@�������/��Iq;��6����kc�ݍSb���|���(��]v.ӄP��|��2pZ�bBn.q��{)���iH�U//>�3z�����q�bھ�?-#I�Nv�i���$*����[a3��k]��D�Z��[�J�G4j�������P�ƙ`�I���S;:�*�Z�|3���}�O�������B�O&1��%K:�V���0�%N���?F�Ph��j��]g��d-�.�1��[��H�)�W"Kc���3Զ@�5�h,�٫�r��V�3��c���������;�Ic)��_�� hkљ"�1*�4���b4.7��Eh�_����	���dZ��[0���VX�{�^�\,���̢,�޾��Q�g��5�{�̦�>����jx��˓}u|�yg�a��d���̽�2M���m%A̎����f��N,BkYO���a����9�J�9kk����z��<~YKh��C�|�no��LnӬ���C���>�Qx!�y	C\9��x��6Jo�!(L�pj�D������ �%��Ի��\�q��j�K���^��F?T��F;�كP�+/�U(��.+E��[)��œ�A�欱���8k��^}�^z �)�sk(;/"8�R�sLф�.��@-?�#�wMjm���(Ity/�
C"pf�ޗ��c,n�������5�����j�W��@A�����A~�����g�8t}q��f)A�2I:+�tBD���Y���{�W�L��玐'E���GD�Du����8U�5�Y��D$#�����H����x,L���Ν�2�v� 79���'�)����cvp�a�>�
�|� ��YM|��Kꆓ��S�1$��4��XSyѿf�lIIbaː��> 6�{�χh_�:�S��$���~��ۢ�Z
�3	�0p��|��.|,l9�ѕ��=����i��������S�A�W�j?����W�ؕG8ԥ��~��o��0XOB����s�>����7�Y�8�	o�Ϥ0f[�~�	����5��R̅�pl���	�phZ�jz�J�F��
�\rҭ�T(�� ' t�v32Bu��G�Pa$P]8�U���j�*s$BR��[	�q	�?]
�g)8|^��m�:x3�'��,�5=T��0גi����y�l2��ɢ���R_�:��a~+_E+I`���_����׊��/\n#�PjX@����N�yZp(AGa�E�&����1�8@�!�)�X��S�����u�ʞ\�Q�tܾ�柱�h�2'+�܃����Lf9	�#��=ڨv��'�pZ���'ق=���\_�$k)'��9
���W�K�<�*U�1��gh����3��4�r���j�S�K3���	r�c�H��;����n�W��ͫT���h����	t�؛��0-{߂�̟DԎ�}���w��\ٵ����:����)��5�{�7����i���Ԛ��s��#��F��y�ݹ|>&��	�-���Μ����d�-���\v��R��&��Q�hr`td�܁ >(���#pU ��W�zP&kZМ���<�C9\��Y�94�2�87�G%�1'�� ����V�c#��W6�B.���0�=!~�]�)��>m
ߌm�C	��O�ǩ�w�϶���BOh���"����3��K&�Ң�ޟ<�z-5��'WVC������d�E���
A-�&�Jrޓ�!�"\YU�ɾ�͹�KgR���6�q���H�ԢPX�5��;�@C����~d���Y�սI�� 
�j�]r�z0M��r¤z��k�_\�j�v�^%��گ�����M�2z��.Y�RT�VQ��*�t��?�_����WP{��$��l�F����]�PY3�����W�>n��g�]�֏R՗@0f����@�Ҹ�35����q{�q T�����_��Z=����	��O����KM�k�*S�_��`�:���lwZ �E;1��O"��騩��YŪ�˺�Y0�fag0��|i��\)��JD�]�dp��ªMd��T$:;6�ۇ�]@�R��LRR���h	�3|mъv����S�,���� @�Q�����.�$P/��@T=�q�������UCy<��.�C��YHn֔'8�0r��}�V/>�����*zq2�U����+A��r~����ט
_��w���m!|�7���>(O�%km���+��q����0 �ͽ��_RK�I�/?�Ӿb҆��\6^����\H�������� 淮�D���V�~�Ƣ�a�r;S؝�I���H�<����ܑ�f���!���aQ֝�@Ή��4����Qi`t͡���i|G7],�2�e��'�k9�*�.�ty]Uǫ�sv~"YD�x���:�%�O�X�o�ɡ��*	�НF�h�Ig̈́	���@8����0mw��Q�"�S��B^w����_{�H�ak{���Rpr�������H���k0��\���~��pk�*�4���0����{v�hRR�[D3�e�
9~���[�G�T�Y�,�%l���L`٪�&F��L2�`�fB���Y��$�ڷY�xv�$��h>Na�Eg��|/�ү�\�Z�g#���e?�#U���A�n��I���;�o����v�a��s���T�Z>�'֍t����V�����v�@<Et���p��)W���e�~l\B)G]��,��1R�Ӄ��Y��_.+}+D��(_Dd�d�����+A��pwZ�����B>E��]Oq�&�@�Ι=����tG�^��˥�
�F�a�O<,���"�ˣwe��A��r@�4�X6����5����P��G�̧�8�g�WJ��v��{�u.I��l��,ƛG�Խs�/n��o%�Is����T�"AZ��">�M�����Y�߯��n�����m.��T���Z���Ks��nC	%f�Y�(0y�)<4+���R�����p��!���9�>h�J�W#��Y�N���[F��Y{��K2��ӷ-��28H�R��ݎ��Tlm������q�)��g����u3~D3��{�Ǌ
-^��t."�(0�p��|��E���(k6�]��M��Sg�Qd��+�ƛ��G��i߫J��bv��N�W?�(@�e]�ܖ�ޛ`qBTm��1zܚ�&��/��@}�N�9_����<P�5��س�E4�B�Ut��<���_QF�9�!Ϥ���PʳDȣ�\ڽ��t٥�ՙ礌���d�~�D���W�03��@�G��^f�%��ѱɍ�,/�LAzT�OO�0�	T�Uc��s&�vEp1�w(9�u��g'���7��g�	���]��e_��?�V��`��� T )!�]�ʣ���f퉑W���z�Nlz!6>3�eb�\�sW�I����g>�|�(�J/��[���iZ.��D�K.���G�����l���IҾ����48�AN��K$r���ɮ�$�+�O��f�����}�Z���^t2,�Z��� ��:,��f��o����}+�j��CA-ppg�	T��e�W�%�����wf���x� c��[��q"�A����(��a�B>�TKnVZ�#(?��q�>0��4����6� [�;b�oY�E&�q?��3־�H�Z��9 D��[�q��
�����d
5��̀�����Ȟ}����{�+�GwhD�$ejy�F���7rr�%3�r����*��u�`p�f.k����Ż��C�x��y�a���7�Th��G&=�:S�M ���/T�1W�>6�����-2J������#��5Iĳ*Ȇ�=�����x��u�-���D��� �|���ś�[��'u�O�!���M��J�)��&>�u�0ȅ����
[��^���簆 ͘��~������XCn��ng�<���P�� +�a��l�*�D�>���|f_�@�.`�*U�'��w'SD�@�QD1�<#�<1��5�]���0����uO�tz��'��D��v�}�;z��r�ǭn1�z�W��ڳ/~�{~����s�^BznW���_����+������$K5�8	�zd#�Ʈ9Hd�f��g��YZ�I�c��x���.I��x:K�V�+eF����N���j�9���B[s~���8���9��ɖ5$�֣t������Ü�)~Zρ����En�L���U�7k�
�)a���A�Zh�}h����E)��R���.�p`����{����v�#��-�X(����0�QJv�����N�n �� j�T�v�3�y׏�I�ΥvN����L0������4E�$l�A��e�Y�PifK���2E�_A^h��OL�X5��Цcj����U�7b�|�b:��J�6�Z��I�h`�'��8��J��ɷS`�p�ٌ�ڍ�� J���p�s
�6
�Kv;ǷP��AKha��G#�9��Y���E\�q�n�@#d�$I���)-�D�	�״�.Q2�v�����
�ʪ�f΁?���h5�u��m��a��q�!y����P^����q�ɒP��% �6聛����YH��J��&i=P���%�c[�U^�?���|�C�6��&Rg�ghP���EA:��FN�S�ɵB�=tt,/���iݚ����í���x�A��|�3�u�VO������B��<s,�$�jSD+b���i!vb|�|L�x>ĉ��8X� +oO)���~7j��krl��KN��?<�O�r4R��3�0��#90(	��/�i�d��W�`�5=�p?�bG���L��=�����H7�u�,o�<A� h!��Z
��=���������R�V��H�c?\�
�F,h�r�r}��������px����rk�|�ϒ��J�_YrD����	l�G4io�e�0�����+�:0�5ЏshMi;�f a��Z����Z8�N#"�$��}��B�/|�Չ�m��]W��?���9|7Z�s�؀�QF���:��0q62������bk{Fs㡫�Ӓxy-/�w�j����P�φ/�4�ZH���k�,�k6�f��Oï�C�������޶��:\Ms��1t�a��À_�tq]��1��;���Dї`�������g:!�3�}O挐��3r�<�o�M]�{+���2z0g�Gk	����7��~���i�4R�mS���{�A�E/��5WBџq�wb����O"Wb?��F?��f�ʻUd��W���ӛ<d�����EQ-�v:+�C�%.o�I�q ���`H.Y�1G"����9,��4�s`�o֡4y%!a�)�ܼ����(2^��k^����p��
Rk<33�턾p��5,Z����c�f��Uq��dZt߃���p)��+��o(����Z�����z4��k�ۇ�2�m�u�.��Ť�R�E��'ja��Icʲ�ֲ0����Bu��!�$�L<0yT���'�#��Ov�B��"�^�y�6ă製=C
J�LM��2��@��u�^�B��0B� �05u��a!�S�n8j*�+	�������/�:�Ǧl�nT��@�97��F������O�
�ob#y�
����P*�8�E�̏F�n������^���
����)�G?T�H����Q�3L�2k��Pw�&��g={�$)_�l��e(�?�*��`s��;���ͽ��DoY�IoO�>�)�5賓0*8ٮ_Mg�����ձ��A���	��n�Jj�$4w�
��M#,l�!���G��3����r�oI��WU6�+��<�?X��?�$s�U���q�-ܮ��l�u��%W�l��
���Ç&R��~^��E
���sS����h
��W~z џ�O{��Q�e���W�N�[��I���8�I�)�� �yVW�o}9�GAJٗ'.�{S+��.?���7�S4T����6�{AK^��K���[�>���	Qw%t6��f�t�SjJ��G�v_���)Lq�S�h~���,+���&'���F �<���`:�}#`��V<޸2a�a~��g�P�2�bmB<��e5���#���f���	��@��4	y1@��B>;�BU`Qmc���|��m�1�}��󧡇QY�֛�:�_�d#�s��¯1�����+�?K���Ui�i���^�+��&�v���s�v�a�Gl�ΆA�I�[�]� ���>�c?t���������۪G�t�����e?��vE�>��ɬ^=�S?pV�t�ErYw��M�B���ފ �����R��n�����8@Hq�t��!�����N P��L6	��k,�_�6��,k�[���[����'�#���c��AS]-}!�§28pF,,T�2(��������h!/��iS �Ь@r�>f�߸�M~6��޹�� ���*��uT�a����~�#wl�����X��C��G~�LUq}�M�Q��&��/[��7��aSEib��Q��
#ݥ)2��>��z�3���B_��CK�$;��p�+@/����a����>^��D���_�c���ԑ��Gm������4�3%������o2�w�u惼���,g�0I��?0K�� �W _�&P�l�����|�E�Œ��YOd�i�	V5��p��h��D�|����R&Ź�~�p��,�PN�mq.2D�9Ɇzb�~C�s�v�,������䕖<��<�[�ޑ����]>h�Y�C�{�l�Q21h�ŅGA}�q�]������9Aڍ��GMX���F �5�@��6�?>�3>Q� D�*T��a�S��*pJ�D|��p�@z�O+�*(�>o��B�z��M4N֤���Yl��L:P�Zl��3����R?E
)7HW��_������{�<�#?fA�ʿ���Kݵ�̚���-��>�!:��|�;��I^̓QF�
г����R����#4�_�ܦ���{alh<V	��o,�����얋�=!i��#V��a5N��_s����HZ�Us�6� �}�nE��Ƌ��ܢ"�4��<(�7i�&�8v�`]#�s�!,"��@`(��5�7�&�x;\�5�[V��R2�0�myF������t�ۗ�t������l�J�Z�$�w�r�eB����<ܷ�#��v�f�6]$\xQT�4N�?�ZE�s�j{Q�P��L��h8����}}�l���_�-7����l�"t�ݲt���� P7���p~�i��SQ�e�A.ZU閶%�?l�=���'#��D!1����e��Ge�o����{Õivg!���k��^uoh�t��r����Ӟ��L��)9G�:�F�����,F�B�Z�֥�'!ͪj��OB8��Ro��[h�:�}�GX3��£��YS�v�0�?9٠�k�W�2���l��=�|2���I��������0���%�2s����O;N��,�=X�~�#�_~=�
�v(��<�<�'s���af}�}�I�K��f[�٢�ö��{��m���~~-h8FŃ���	����<\&x�&�^��A-�S��5�6^�mM�ِ��4 ���Y��o,���U��>ϝ��-���1��j�Z�8��A��/xQ$7\M�1�T�����F�o��Y���F^�L�D?����k/W�}�C!Z�V���Y)�*�N�iP�d	��d^	.D�a��#�s��^o�"��A��l� �j��ӵfHh���A���]����3��Q�`6F 1=�9��=� ����lQ�������]��.9T��!�"���O6���{vN�}�9m�GJS�H��aFs�bh�nz��|���Vn`+W�{�3ofb��_T'� ����.v�'N�D�`P�2�,\��ӎ �Ņw�w���D��t��h�G�v�V�Ԋ�d�U�R�se����g.��T���E��;?�lg�d�x�!9�[�@e�t�DٗC�"|����&�}x�+@���ÿu�Y�c�0����%���
��M��Y�`��t��l%�R��QF9Ӧ�dNn��F	����jH���rHX�rT.��EJ6U�.d�IM�@����P�G�!R�\��rb�U�����NiP˺�a>oޅ5u��j4��nI���T/���mmB�=��?X۲�d`�C2�m���5��Uoq� �ь��X��o����Vͩ��� K�2�`(��s�Iz������_�S=�S��T�]H�$ �O,���R���5��;���mf�> ��[]���Cߎ�3mΪiz� ��$�nR o^B9)G�(�i�����v�Re�.�	�0�����da���*��U�߳����J��ʋ4Odػ�B��d���}&�8�-��~����AN�����[oJ�#9E����;2���X�-��K�caE���N���t9Ύ/N��Cz7�݂zhG3ܫ�r�ae$�fF���,�V��H5i��Pk"E*y��-��)з�m��B�"-�w8���]����q�U?K;�S�i�S�~z� ��"H�+�
:7�0�Y�@���3��#~�F.|�J�M��̷a����'�A�N��2�'�B�����/�-�nIؼ�'��6`�X+Ҿ5����@��Egr�ġ���I~,�`Y����S[N�N�y+�(�J�avq楌}Zk<gH5�N/9zn`���f�Z�T�t�|�����j�ʅ$'J~ �h2�J���d),��λ�U�����H>��f�{�#C�#7�R^���!%�S�%?n�����&�`}},�A����ݫ��Q0���Z�4�V�[r���{A<�BC�4L�ag�}Lg�ÀHB!�=52�И�\��w������F�A��2χ%�8B�K�'��g��l�L��o=�ňnA���ιUqݹl͉CUF��
��p˰(Q1�&��6���X���wmuHo��3���؆�XՖ J�ڥ�4���S9Y�;tėZ��"���K�j��O Q>ns�ūt��7��y{5 �g�o-��J����ӝf0�Ś� {qw˅�F�|N��!�s3���ю�Ϙ���_���M�@��Ք�[p���n��-pi��u����˟��֮c��dcv�ɿ��*R(��Ϊ�ɘ^5?�l6$�DΥ��I��o�;�,�G�{+Ĝ�'?z��i����݂� ��i�y��W���=NB���,�����Тo�S��Fγ��u_�V;���X�m"_�{X�����RSizP � �������f9�򇢕�Z�OA��i@��=�_%�̱ۓ_;4Ţ����z�����8��&ذ["0�x��O7�.��и�����̐�+j���a���2&�ȳ�l�8���תR�/�	�δ$�z�����}@�a��2�«ᒘ�R���`lL&#K�a~]���k�;X�^�g�K]���1=�3#�*�4-מ��O����x�|nT�6-����?IcDE�>�O�#�����R�kdU�#|�W��v�!}��e�BF��ұ)aWx�G:�e�_P'V��}uװ..�Y��3P���B�%!��L=�읦W<�����6�{)���&���i�H�FdEK�9;>	��m�z��[�e��A�I���l;{|��o��3�uj`JA�Z|@S�#&��s"`V=��0u��,����_�k�b(��u�I�R~��B�ĭ��q+�E�A!��8?@����r������S̢��¶����^<�����JM���[��n�.m���'�5�k�sU�V��ډt�����}nĀQ��_1��f��~�<w��XZ7-I%F�Y�a-�B��κS�=&�y�'r,��O�x1���8ˎ6��;(e���y�R��geT�@�S��4�P0SWUK�1�Ҽ59�'��І�Bj`�S��o�98z�����&	�b�T�I�]���6]����}���<��>�s֩����!+o*�:3��$���G���ۏ�(��7�yM���DVקh5�w�7y�+;l�G��n�x��p���1ޡ;�3�9��<ֻ���o��OsC}){H�В;F�)���Ϯ�h��rp���GI�b
����O�Y�+kV�H�y�����i�0�#d��F
R��bŹ	��K"r>����HR���}�o)�����h�*}~E��淃Z��vq1�Ǒ��ɧ	�$�Rwk2=g��c+��\�<i��x
h��� %p�\�5�س��V�d���WC�����-d+]��vC5d+Ʌ�\n{��҆��'�:���,�)���ϥ����ж۷�
��N0����a�n�{d[	�z���l&Ց��:��X�z;�`��f	 s�Aޢ�T�aK
�����w�9����Ŕ 5�+x�y��W��e%�)�+���M`��ߨ�K���\�g�L�<[��`p�1�u��s�<���޾D4�5  xcno�
�X�[����drΈ�W��%mo[��f$e�����+�֏�h���H˕�951�4.��W�C�:�d(�� ����3R�O���a�yȔ�s#���ğ��ǋ�4�cxp
�,��Nع7"��~I �×��K���=,,���o��Lm��&��qK�f�{�!�?�ۥNx�C�S�ٓ<����^Y��g�&��mS���o\O��"�Ğ������	,���2J�Җ��ve�n�٩����"��=�;����ؕ ���3]���u�37;/��H1e6줬A�]�2=�o���S�S�$? �?T��6KV-�ۈ��������D+����z^a�ƌ��D_�5�oӨ�������;������@p;��%�$RPɍ��`���FhT�M]������Z�܅��dD��~�/�t��кu��ISD�/��b5"§"N�ӰښF��O4��H�J��fP �g�O�︂aH :��c��"#�:V���<0�����Օ��p��ė��g�4N?�_�������F�7i� fm�3�4���XC0*�j��̻?�)�6��h����k8]��E�Y��,d� �9r�E|�d��U�7�F�i�XKG���.�J�o�c)T]ɷ���Z��=������*��cKD�1��4��5�mQ�X����e�Z����B��]�á~���RZmC���g4��f,6e]�b�1P5cl[�k�:{ ���Y��R��
��)O��񗪁�!� ����)�Ps:�7�2w��l�G @�k��P�\'hK�s��Ӑe�����Z��.���ĿD�d=ŅV��'I딭��n��a�`C�N� �'E�?ީ�/�28j�a�Z1��M���veܴ��5�<n�Ͻ�Q��ٯA��|9k.qIa�C��$�/� �����ݕ�H�T.s]wM�6>U�y�MC�ڔ$�;ST���@�>�+�,abm�#��G��ג@����}D�%�<�S2�kP�4@��m�^�h��G��8?�$�{�?��J���q����=
,�a�r�]i�xb��O��F���a8�t�E7�TI��̸NN�}Vm�D��x㫖+1��g��']�p�,?�&���=�'x���h��tZ��+���5�G�:dy�a1�g)��3	^�|��S��H�/���@C�Ti�iI���ҦT�jg.����D�Pt��(	6���Pk�Ƣ���oi�_����B��e�M��,�N��+k=�f�}%�g�>�A>V���7��E�Ծ����A�<��W��=J�¬�a�)L��n�@�(^z����>R�����tn�.ȷ0��p��<;�� Pb۲7`�q�!�w�W��*�&Ip������Q:�9�3»��q�!����^�|M��&�;��P�����[��=�]J�w�v<|6�6�#i���j���#Z��
�/��ǩ��M�>�l+��ֱ�o$ی�X;���u����C�Z� w����Y�W&�!�8����?u�)��Y� I\D�pB_��E�1�;䥈�������l�QCuDO_rq����#
��d�����B����y�"��o�}AN�&4���;�7j6o)%6�&�\=2f��z�;6kP7�@�-8c�����W����eu9T�ԌXZA�U=Ҭ?��UK�Ŷ�~���t�hk���?g�=���"fGR����1���J��¶� ��2b�p��OV���^��ƌ�����;�wB����]u��ͫ�K5� "iSB,M��v0��.��ku��O>��ɶש��ٌbxiD�-�M�MW4�W��j���M�5x�&�51B�^�w����/�y�$D�샃�T��e�<o�.�I�A����M�DC`խ���� ־��9�c�j��s��k�v�:�.��4�H��>_��Ʒ;7���G؂oڟ����F�2�W�@'hN}"�߁��9�<��I�ħ����-H��R��"��'���N�E��K����"C���<���������Ǫ��BO��8�=^�o<b�O�A:!uP���qL�$Wq��DH遙�#Fɜx��6�Ԉ�D��I9t����5>@)��Z�������E�P�h1����"޷����<���vk�+�j�^����}؛"�bM�Jל��g�$g��e|s ��c��	�-Hx�W>��ߘ�x�æ�2��:vTî��R�#w��c�$.Wh���W��_/�Ki[��*��Z���헶�m��y�82ǂR�7ZJ�l�D`:-]�ӻ��t�蕷�X�]�h������Β�����74����v=��$���-����(N��3��w_t�ȟL��0�T�B)�S+1R���?�z���1��L���:�Z��a�?v��s�0οQy���)x-��T�M�il?����[��:r�ʘ��/lcm��y����]I^-�N�/��ŧ74pkQ��_�e�g���ҡf��%���]F����̭w��|��"�Ui��e��J������,Q���}oR�L���C���΋�y�����j���y	d���Xmv��&(�T<p��'0����H��ܙ�!´j�q��!f>J�Jp���U�,,h��UD۹�% ��T&�p����bU�O��ɮ�1l���}�B��g]��Ź�sjʵ(O�$�yʃ����\�K+@g���Ìq��OE!��\��W��?���N5����a^�����X�N���y��-���=_H�&�-a���9[X[��<�q�mO?�D!�+pZ
9~�TQmʗl��)H�����R���´���`�B��7��N�ab�y8o^1�&D�2�y����������r9Xj�}~Yl
����}L1��'@�N�O;�M��D��R���S��0mt�l�_ A��ğ��}@�-TqKX��;��I;�=���7�y)�u�[|���֦��.�°2�L��)~}M�"Ë��Z������{��$y)R��okڴo��Be23V�n���qȩ�,ɴVMfdV^�똊D����r˖I�ſ����q��lq�'*".�+4�(���#�m��W��2��^x$�ڢ���IU�\��R��Z1����ϕ�-,�m-02'�6e�PB�%��#*6�Ŭ�9�>�8˕:�:EY.��*גTUR.B���a�C�j��1��Hs� �G��T��v�ȃ���R�x �g��=�	�x�E� �#MzK��it+,��3�rӀwU�G���Bz&�6_ŇU��9S��r���v)��#-��"���(��!�[�Ngڇ��t捩��F�NǟP-���01-A:�<-%�7k$`��6s������2礑Y�����>�(�a"��Pי�W6>:'b��v5^��d�΂�D*GJ��T_[iX[��|tr��m�n��<+�(Vg��@�Эۆ�)�B��F�8�ֺ��g���2L���^���`�e t�PRX��&�%M��4D�����.��P���Z�1��i�	�m�A,��"���WH��3(a:��N�;�v�;�zS��		H�[�+� X^�d�^/�_�ۄ�I-�����kIϹz����ܕ���G�A���q�~�.���|L�|�@�5X�TԵ�������(���	� �����`@��(�T�/�;�h'�Mj?���8��`�a����¨E�ݶ��Tu)GX�fkS������Uk�u��\V��z�e��%T�^� �4ܫ�Z
�W!����Ł���hgD'.�A�R��l��\�/y#w���5��)a}E {D3�/`6�݀������C�7�{���[�0K���+4��7$9q�F�iz1�q���`T^x��̀������h,���l�
�L�L?V�nb�օ,������NZ����t����ZDr�0��K��%5��D��/U�ی71׬*�;�w������l���j��r���\�N`i�`��=S$>��;=jT �1�%�w4�F��0�[�R��=h��4akLO'��;_�f��#��c�+.c�?a1cC�EU�V0�FK4��o�QEh����iL&�ڥ���y|�����IN2`�f4A3O���<�o7���2�ҹ�r	���1C��jǶ���p]+xc��}�l��2.�P�ܖ�P��?"B���䟙/j
���ϩ�Ѣ�������' 2����nso?=<��BI �՝]g9~S�����%Va��E~���}�¦B�J����:+sӝD�k�`�K
�+���Y����N]ãU��Xh�!	�E�Y�px�%u�^'$�2��x�-k�5C,�Q-q:�7 I1T[!�_c6�e�Hz�!�U��U������N��q�(rl�zY��e�{85
��W(T� ��KWeP�}CU�h_� ���_�_�O�o�P4&��>�Vo�������x�	B��M����i6֊��+�Td	Fљh�%��)3��`	�Ep
���Y߅6��=���&神����������z���
龛jZx�4J��>��+@����	��ԫ�� �3�ko��˛�����&t�%eט�-���׺��dEO^���S-p�&a�9�|e#��$$ �7��+ch�����Peٷ�B���X닀 _?���m�ߏ�ڙ����h'��}X�8K5]R|�Y�"�n��"����P�>�Jp��B`W���ƽ�$f���I�:N6�����TAev}�GW���k���Fä_m7� ���d���h��౻��d_�ėgu>��ӣM�:�틈�Z�$�\� ���]�ran�άUá*fT���C��D#�W+P�'���su���vl��b����-#�zC����M#�p���{��M����������}`�pK�$
Wv
�4t��k��Yv�1���=�QG�����x�2�z�/]�0��Z�� ��{�BT��a�I���T�1�:9��1�Uv#�%����*˅57\�>��'kߍO����SV��
�j-�[�z��Ә�YR�R&r�\2�fT7��(�a舫�kS>(uV�S��
˨�UnD�x�"/e��ä��F�5���p�`1���}J��M���?�}���O�f�wԮ�����2*���+��l���φC�,[���%�
��	�!�VT7sۺH���;ľ��kCEA"O����-<Ż��CE��-��+�V�z���ZKz���#�e�M*Û�5'"�E�������֎��у��V7�,抍P /C֚�4L�>buW�ϳlq�H�ˀ�//����}�@���]�L��͐� �7	�<��K��,�S�f�:����(���p��O��r�L�oW?u�ݶq��T+(��N�`!e ����>��O֏��!Qs
�7��s\e� �$�w�)7e�K�	v
>\��5�->��<�qӓ�̡���$�������K�f=���Y�*u�"���<�G���{�*Z
���i�]��Ƕ\Ue��8�I��@���t���ogk�mŦ��5��B�M@�mG3�vzzK��u�C�\\���lk*�ʹ��g���C���㩕]�f�U-�?u-�:���XKq*F5Wi�����"p&�̿&`�2��?[�۠��~_�ނ^�E��P��fRu���Á���I� ��v�>�Y及1���u#�v: ��
��h�6���b��� �ְ�3v�A~-�y�C3'Rg�z^ ǲV���f�^�[�QCML��3�E��V���e��i|��جƻI�/��^�me�s�n�P>o���s��3Raу�����~i��B�C�G�4����M�f�c�>����@<V������/:)�Sг�M���F�U�m	j�X���G�mW��X%/�MŔaKWX�ԩ�W�l
5�$��CeF���]cG:�r�I�%��xM��1̳	��ԭkGȦ�3B�v�-=�u�������i{˅fn<�U7����!֍2����Sy�_�m�$:��@�U3�rpP�oIF��|�$�W�7¸?tH����m���ץ��U�a��'�o�ˀ���S!�x����A%��Qv=��n����%���;�e�8�������&�>X��l)D�~=|��Uim��]��*��\�zp���/.jy7Ɉe�wz�/�����s�j�Y:�e#Z8�&S�=�)��r���_6j~��{?����l����>��>������)L��c�qǐNً#pI�,ɏy/���,��cN.+P�?A���w}�Ӌ	�{��p�Ƹ�Cc���^L*�o*Z֡�?�h/�����ʖ��)F�����t~���4�`9�;�&�]Ђ�iU���%{= �=	�V�>�½M�H�- 7��4U"�p�zޗ%�'q�q5_>�.?:@�������#F���U�Z���ȫ;�K�TP2��o:�������wG#)X�5����+6��������
u����!ɗ,@��>^!����Hk�-��)��;���N��Sw�"0��������Ԃ������b���3P�e!��ڬ������Ѕl��_㉀���fAI���fV��=���N:ʆ���[z��P���ق*%����$��17�P=������s��{��"������;���PVV���̓\ۃcΐ��B�!�j�pO˫X�S��d���k{��CpVveĔ|@��E(������(�O��Lb
�����.��,�T�P< ���Zf�����I�c�4'��(�`��.\_I����6�Ufd v�ޟ�.�љhͲP�>ڼ�*,�)#.�
��]�zP#��
�94֙����߾E<	&�0b�}�����/�L��^6_��Jd�X��X���M��fR,�}�L�M�F-�N���blf'�*E�)�E��)zܩ�>����*�n�9���S��{��f:w��V�>�>D�����I.W-�3
�$␦�������Wr���>�k��I�?G�`R����p�K ��{���ؔB��T5��фAZ�e'�s��� [D��	����"@7;I�ja��"e�ʠ<r����M3�����dP�����$��'�rջᴮ�*ԃ��'P/D;��
�I0���Z�l�T���f�������=Iq��g{"�U^5�x� �(���k�r	�l�2~����r�4�"F���l����d`Lks�S� *��X`����~���
��I��Ƅ:�����%xd/�r~�-���� ��x���ď�b�����5w�b�c�:Ū��]*S�y����Ɛ������������v\���1b�)F�7�8������Dj-B�^��z ���d����J2O�3��2\�9!μ��m�׈q��^g�J֊p"
�O�Qѐ2@�S��Lp�s8я�MAD-K�u���3���ׇZG%�%����cмTLXH��\<�c.\�ns�C��|a |�n�X�n�g�&(��݊gq�Bb5O/�:���� �����y��u��W���lMb��JRe����b�k����W��y�.����A'm��6g|F۳�5�Y�'_����PGQ������58W�`{���{���5FE�޹]$�v*�sz�����;�E������Rs�I���j��L���t�m�s����)��O�^�t��/�&�>)��z�4$f�^_j��3=��1�(�&k��7�c`ZM�O���(iDv -S%h�h�z�=J�r=�b)�ѰV�o�t*Y���u���.���%��R�q��ꕿ$i�`�B* ���-�ܜ5�`b�c��{k0h�2�}�&��9�_�Q��d�A�*@z���ZD_1D1��������9����E����b�d��P/
�
�h�w��j�[���4Ze�_!!	�E匿��%z�������e�Z����O�![J�A�22��`�<|�! ����˟m�\�J�G%즆��]fs��xrf���
�٭�2� ~��ڶJ-l�� X�;,�'�~�6�>'Q��ٜ�/�Q�y����1����n��|�ќ����/���t�K���`O7兏�O�c�7��9�SlFD^<Xs"��wk�$�F�\��k��=���������,���L���@�*�O?��v_��_Hő|��>��e����r��ǁ�} �E����`>���բ�2s�AW�P�1C���`Rc 4��o)|1o<�9Z�p��KlpAt�� Y���Ծ��vw�&�m�L���`�a
��b"�)Xj�<$�s]Sy�J�%�kP�]뻬��.Q�����d�9�Ђ�R0[8�-��ӏ.��"���3j���^��Yrʾ{p�'[ȑX$��+�X���`�n3mU\!�Ҁ��[;51�O="ΈEqRw�б m�1��QÄ��"r�L�f��#��{���/R�1����d��"C��%Fo��#��J؏z�*�9��qX������M�_X�,�aKxU�y�#��Z����ą EhJ��[�����0B��PW�7n���[�,���XZJͮ���ݜ�q%�晓,��sr���?��AA�xȡ�~�����;+0N��8���9#�M�V- �EV�T7�ڷ�����4�)�1�	�D6ޥ�E�ީ�*��ͤ\���Ż���4��i�r��d7Q�wmC�����3�W}�Җ�nq%J�+0�(W/�A�(�M�
�H����[8�<�K���އ�&m���;ֽ$�m���(����EB �������u�ϲ��piV�jɗ&1�w��*ۮ@��2J@C&�`��ˁ����	Y�g���6���Fؼ;s-�����tOf��L�V�Yn�S��%�w���.�xW��S���_��<+�E����5��'U�Q;��f�8Ox�ʕ-s��"#�x������hԊ� Z�5U�y{v����j% g+��|�H�<�tU����*���dӂ�r}ѐ"�Vc|�ȃ?dg5�{gI>ɊPtR?ݏ����	�X�ќRy^AD�L}�,�b&�y�eזpC��m(��>~��%_�L|:�wֈ�z���K�sk��p��eICJ��f��v����7���xt"4�MkE���V,���XVZ߹k�����x(.���乗�%�^�R�����å�-�M���h�0}��r�d��
������	'��v\N��4G*�+�q{�6S�����7S�?��79�?L�h��zL��2F+�m:�'��^�����c���2��-E%)��D��1'؈[_�����Ƙ���P�-Ԗ�9��c�� ���*��?r���� *�}����|c�U�1��eֽ�w���ilTxKH�x;�v0b�}�au
����W���{���hcuRFߘ���[��	����1_�T�szl�X�T�`��z�PR�yG��L��ٟ�	�`������l4qX�kPFc�����r8��H��(���9uP@y%�Fa��"^g=�D4).�q^D�ܭimKڱ����Y9��Fy8����ث?WfKWD8���$��M�,��]���cb���\g��j�[VX�ֱ��&k"��G��+��ǖ�P찳X;��Q�X���,#��Gky{�Nå�l�����΅��^�FZ�Z�1��` z�;�n��?���B ��ɝ�����Y{�褑l�?�C��ƚm��#�U����bJ����"�QTi2[�W���"�#�@����F�g���W� �����cڂ.��z��t���I�+� uQ@�{=�l�0%U�^V��n�<���\���恀~�fS����ZH�^�8`V{�ax�ƹU�+6ȳI��rU'�	|�f߮��kÆe^��q@WC@Y'|Ov�늪yWm�5������No�B:���Kw��ǢJ�|���}�T2�E@���3�GBF�X�����T��d}\�&�S����|ҳt�k���iͽ��M�B�	z`����i_.����I��gV����f��
�<��-9G�u��^�R��Y����i�n[v��Ep��	�V��{\�2�d�A=i����R�,�9�Y�����M�����ۤ:���v�C�;�4�)�%�*���PeL�}-�x����(���fh�I�CAMZ��~J��WA����W����E�t��Y3_S;JԖ_��mqE� �S��-��a^�HYv��/L�1$͆�iӱk��z�]=���S��B�����ǻ�0Q��a�R5�%�S�]b
r���8@8��c�*Z��*���^���p�X�v.m4��C������*���g�m�!
�mif^"�	�7����~�X�C����R)�wV*�gmd�t���姣�n��p:o�)��ׯ�3ز�$L�9�`����t�+�� ;�W��=�q�vظ��*4ތU|�Ԫ��W����C�A�T��D�;>��˩M���]4��@�mj,���DC�����'�������Ho�ŘS�س;�v6+��R��of���0b�{)��愧�y��Q�L���%'��8E��uX�|��%?��~y8��	�@)4z�QdF���ST���������GI��t�6��%"^1H��c�+�%|�����^t�D9��g�/�[�4v�
L�_��!p��*Z���D���z
��W������β&��/�+M`��w�f���nk������S��}& q��t�<����h��p,��U�^&�Ox��`s��c���<��g��F}�a��4L��)��=/�2)`�X8�s��U�=��8/����jR��?yF�yL�a���MbW�5��������7���}P	K�����G}<
�!g��߁�xa�~��S��OSF��@j�v��S�ؗ����r���,��M��ݎ/��VoO����t �r�:�ezնG�'������zs�(�ҀW�N�N�z8�h5��řA��;�l��H�>`�6���ކK��ډ����&�]I�%`��bP���O��焤9�2"^�t�Ue�=����)�V�I�����O9��1B�*Д��K-�v׊ڻɑY���[ �.*v�V	�#|��Γ�-
~�H�9\���rAnΪ�'P�6ϟ���On�ν�j��&�`�`�J+\�t�(�=�sGj�X���p#F0.]�JD��f»0�H䐧Ya����]+�b΀.��l��T9�5O���9jh�V��LM7�fI���԰�Z)N_X&�����`N��j\utq͝�/�0<	��~%��v_��J�~��9�bcg��j���=�壿�t��/8}��
�N�lH&Z�$&+�_��_��TФ�r.���r��1>�b~~�I/[r[0x�Ծ�wV�F ����&����\;�Ŵ�3�4L�TY�r�`��<5%|F�?�u�bP�@U���?���ge=j�vÌ۳5l!3	Boh������@��-�M��Hh˥���mʾr��Hu��m�:��1:����(.OX�L)BA43��<��09��j`�y�6�c�FС���� �����H�����$R�x��J8@9��%��i������=7�)��w�Z QM�tz
uX+�B�*?&gNQ��,�ʈ�qk�I���&}���v���d������V��Њ*L�׍@>Oe���1�_U�-<[�f��4�Xv�b.��Ʌ���O��9�U�X���+AT�SvP���2츱�{5���C�����jގ�~.��pT	�̵�V��_NxǤ̰��GJP���kn�͑z�A��c3AZ���x�a3�>�_{�ص_ya柯�^C�Q&h��Z�� �K<u,�,LOHj��ű��dl�����x���_ >�?�+ss�����#<��*�(�T8d��_�u%?�
FH��L���;����L�g%^�B�w��p����
*=
��l�I����|e���>#��'��j���=��9����|܅�x�61�~~`\E��r\L���S`�ID��o��l�}-�e8W.L���0�c�)L��Ru��~u-O�[�X�疕 Q�jHl�+�����Y=B�+�dV��6l��	�q焢�F`������V��ήN.ΰX�/�AG��{�M���d�Kˑ6j#��ۮ�i> 	q��n~iR�l�1E�wG&@#��<)���{��`}���9i~�F�B�`����%�I�R�UJ}����Y�B�i�'*xf@`h)�b��!+�V�2����*2�r�';v.���Ua���B������r�
����]~�e����)
K��JЦ	�� �5��41�B�[|��w)TR?z�)�b��&�cZ��/i��V3G>�
���ޛ���}�����!�?ߧ��r�����	`Хٝ��)��,��!4G���=8�/��b�ʍ�L�om��[{�=?��/oX�C[�H��|���HsS��&�6G757Y�Z%hX n��"In}<a#cW��!2��As|�����3�ﻃ�����^�A�$�B>�%��í��]����m�Ǫ���H[����G;p��7�!�e���H3z��?��W���Չ�2��T���?݂��K�C$��S�[�)3��d�L��Ǉ[J�h�����[(�1Q�^X�q�47�ҨC>�ҋ$���/�1�%����	=σ'r��O��� )�ܹN�*I�hq��$/�'�!.��{u����;F��ؠ��ତ��1�x7� �yR�a��T	ԟ��g��aT�\�K
l�>�đ�@mb�9^�"�WՀ$W�Q�*L���z�{� o�a�ԅG�0�۪N��c,uX9�m�4{��P�d��f?�����*l�vM=��@�!x�o�x��g�UT�E*����b��3 ����� �P�ad���}L��y�@�9n��f4�p��6IqI�W$M�i�B������L~ �X�����=��9��6o��Y&E�j��NOU�t����僛ӧ�����	SlfU1���<�_�80-�^Y�:��[T�7��?��Pj�eL����Y�+�A �
|����T`ŖfL�׏�#I�`j������1=X�s����nM�/g�����Ϣr��>m:���o�23M�c#�jDe�`dTP���vNr�����Kn^!t+�x�x�\Ҽ��,7�mtU�Ж�遌����7L�B��t,`�9c�\�����}�~eY�3�U�Q��\k������O-����U������x!_� �N����j��z��@�[	ƈ�'�WI4�u����װ��J;N��TI轉��͗n�On�N�����F����ZMt�����V����谘c�\��r;���P�D+��<�a;�Z[��~=��x��ij���M�7�w�<�����1]k�c�d�T'Jl^�b9c~u��㏸�'k$��uZ���|W]!�K)$�m,�3�;%cb�A�tB�,�&��I��Q���<e��W�?A��� s���f�B=ǭq�tx�@n�?Y�K�J+w�|#z�g��mQ�1����
w"��!�^�wp'z`�B��J�4�&L=aJrϤ��� |ؽo��2�<��*h��U���dW`i��*��Z����󖅬紊����1p�K��푹�3ϟ-��WM_W~��Xϓ��u��j ہ����!�"�D���Izd���q�h*�`��f�ȼ�]�'��W��σ�QC'��1i���ܲ;���B�[�8 ��@7��eÔB�ǅ݅�����ڶ5>�Ei^aQ���x��(5�B��3Z�����FhO*p}D�!gX�5��#�%�|�l&?7-K�!�L\�4�eF!z��!`��]�`��������Q\��^�H�V�SS���A$���_=<6젭 ���P�u��{�X8DUf��gm��G��U�:Y<N��BB�A!�3rڧ��$�m�o��vW�;��^�QKu.JFV���,�w��(Џ�k�9j�c�iU�N���&6`�o��B B�2?����!1	o���FE�x�h�id`P̈́GS���ζ�ۗ����: ?$ϭĈ*�I�w7z�+?6�#΅�W*X�P�ؚ�c
�@�:.�J��v=3$
5Hլ��^�ػ�Vb� )��%z�V�fS�x�]�\��uU�Ek�R�\�XL��o;-���ҵ%Tt�Z�4d��A�,H��<�%�d�a��p���jo�ɸ�SaZ�B���VC
�YL���zX;��ңC{֘rcF�����Q����@=:���IAB%+��O�i�G����GiXnTs$���Ż�5S^�q0>��~K岊�ohE��%,�F٣��D8BW4�|*�S�T��͜�������3��i�}�ĝR�?���kg�1Sbo�}�	]R��,ݟA��U�%=�k�t�@����KEU�!�.j��m�&(#���S�l�x�
�߄%�{}��d�Qw%0�����	�,Bx�ǜ�v��>�.|��0|�YK�ril���y�e�?��>؇��>��S�YS~����]��|I�/H��v����+���j{�D0��S �պh��`��MMrb2��h�^?�蹙'Q��҇�%x{Pe�Z�>�i#�3/&$(R;aT͟��"�k�=�$�A���P�v�}�_,�UQo4����✉�O��z�C��x��m�>:�Bm<u7�4�#��7���,��g�V��(�~�'���x��.�K�/F�y�	47B����k�\�<+�E
��ld0�b�|.�tlND^�@욁5$p{���?���;�m ������,?.��!]��-�����X�x�?�" R��H�q#�B��烙�@�@Ӥ���Hf}�b3��F�t�q�R3�;���X}':����Կn_'�ͱ5ď�"c���]0��Kq��I!�lS��Z��F	�|�a:�\�U�N8�#Dj�c ,|l�B�������gXՒIQ����\C~���X�N�MD��5��5��EJ�����*	p�E���]��%�\FY4���w%����s��b�dys�86-���/�J�����4�8w�j�^eר^˱��8�k����E0�C֬���� J`��t��p9�nP�s^��Rҍ�ᦋ�Q8
e�l�f�t#1�Q�iW��4� ��2�pg,i�Ζ�H�Y:Y�=8魯�(�;��	R�Mo�6�kL����Fke�[�5ػ������3Z�"�*���5����I�Â�LJ����4��Ű��D<��5@o���E�=�9���߀M�;x<l���1Þ�Wk�������\��:<�ƈ�m@@��aC~(�����B&o���
��V�k�z�I$w�{�Å���ju�)���Y�"�I�W��4A��vZx|��tB����_mh��k+����&ް�E3(�}�� �|_5[2����vߜ�o95PQ���z�G����9ϊ�o�{�8�)����2�}m2�zyQ�m�\��H�mY8as��#��R��k
9��C"�+z���}ViL�%��|ay�R����h�����������{'�F0A�c��F��kN�/1bk��Q��{W����K�G���T.Qw�s�ώ����%ܞ��h���O�2˳2��l��*8S�N^OP����m/汁��;o�a,~x�38\��s9�M���^���I6�����@>dw���[����(N��*5�5ͽ�~����ȃl�x��36\�y~;�QG�W?�P'@Lg`�y�4�Ve�9N
�j��vl�pZ�f]�T=t��w�Aq���|�l�񞨈$�0�T���ѝ��Z?�eY�����`F"P8�i��p)�Y���qW?�+��ґ�����R�D���>��_ڑ�U�p��H/��B.�ދQ
qV������"�����2�r��Ս��n���!H�"�R�g7�)~��������$�ty���I�,C�/]�!�)9��G���N,�@��
E(_����%�k��n�j�U�-����I�^�:c^*9N\�[9��&�ڔ��{|m͠�ts+�/�]����&<�n8YH:Ƶܑ��������iR;�Y��M�I�%	�ad�u�2T5�hcdE�rW���6� {ͮ�7s�o���E��z(/1�?��ӭ(|B�ŏ����+��1��5�9%�1A^�R��i/<�"dl��o�J��h�dAO���V~��L�t��B�i��=�y&,&�s�d��ct�"@B�{���$�$Y��4RpϬ�q��9җĻ+��*Z�� S.�h��[֑�[y����B�#�+]�l΀�L,|�`+e���iMH�a���7R=�	���?����D��:$���mu;h���HA�W����q���;�e�F?<j�8�J���5܂M��8���1��>@���?����x�0=~���1j�8��5������o�
4����X2���c�����Y�+����>F�S"7�	�L�EQ�WJä�~���^(�};����o�K��wq��rr�(�
4D�
��ŔKTb��d&�n6�o�hb�)��>$�vr@�9�G��'!F�)f�B��%�R��������������֍��3)t��}Ţ�ZM���L�XBV��-�/H~�af�33,�� -���0i�R����ɆNj{g��x[
��rl��@��1�rR��6� �lyݽ���;�����3(8��Sk)�h:����G~�u����P{����~�ݾx���W��|t�sH�[��Q����F2}�# /���
Y_h]�5����n�k�V�*S*����.T�LϬo�ǧ��bW�ц�˯o�S�JQ�J�R&H~�Z:~*�|�_�
�eY�d���P���� �w����i�cP�����k!/�iv��F����0�fls�u]�g�ӭ�k����^~���xj>n5�lvy��o&1WA^���t��	�qo��j�ܑ;���B��#C��d��������	b@�m��Pf�~S2�N\odؓ*m����@����FOih+�ѫ̏[T�����Fҥ���8����t�A>��@�<em	n�6Ǧd 9����7J�7�Q�nq��^��YW^7��-5�YX	�eK��'�#u�,@
��v'{�o�h�<�pO�+�'���4��<_ X÷���[��T ��4�,H�G�⠴/[����r����FDg"�'G����h�
�N������x����3�A�����]/�^�!{[���(J6%�&)ս�[���Fo�88a�P��\|���K
{��)_��\�]�|y�>�Q2��f#�5�1�׷h�L.B��M�B���S�7��^�m��1�uh�wT�B����տ�eP��7�r�K�x����`�Z��cT�]���暱6�A+0�J�D\�z�?��Q˄uo/\RY\aq�\J	sY���#Na���}�MH���1-{��C^g�`��	|�4�b����	W�9�S��#��Rؖ����/+�|�-�j�+�͡����,���aA�(Y��(ѿa���:l'�,��CGZ�N��NN��Lյ�b����sjp��]|�ɀ<#���-Q
F� �J܋h��6�{-��wP(�ʘ/h7���;����wU���mk�t9Sa�ݛf&)��.�9k�d�M�w%����B��&��_��<��X��Ch|�n�B��Q����uw`Z}�ں�;mk?���:�1�$�|�uZ޼��P�$$n%s�Bj�0�(�X
yF���M��p��>�2���U�$^.�g̫qH\+��?�T$w�QF�יl�>���/E��!��Z+��~j^:i>/��K�_�@ǔ�.�j�p7�o!{;�� �����p����Ť�o����v�B���\3�.��8g�<�G'��rU�c5q+yA��Ƚtp���|(�s/�Q��+��K��g�l+*;&�� 8��&g�w�k-��b�\q~����8T�	5�C�X@
��3u����n�߳�C�_?���}�D���q֛1�p�P���]����F��ܯ�Q�
yH�xx�ՙp��	�;�x��4��s�gt�jF���-�ٟ��@ʤ�r��P}�W��k�#\�:�`��9��w;ЊSF��\%�j��
��$\��\�G��ia��^�����Lm���뙪�����TޝQ`�L:�� k�0����(�d�!հM���ZL�l�
�ݩ0l��S��D㝡d"NL�(�����#�fᏏ�0T��2c�����{���*n��"�c����L�5�� ��"�S�ug}6*��w�ep�1�=�j�&�X�`��a7��2@.�r�n�`�� 7X�6�8=��rm�m�u��*�캹��ՠ�ί�$>A�)^��Q8|Zm�2�cC�J��`���[����S.ȉސ!0���s�����!�����,�8N�:�R�Ct(t�S��v�XJ�O�F�>-.:!fkF���/!�c�����
�u���,N�����Ń'�*��P�8�{������9{7r���y!�}bpɠ�1��ZΎ�X9�'��q9ܒ}}E��x]�ǡ���p��$�
-"�*6[��������壣���/����:e2�X�r�C17y.��X1���8��F^�%nЎ�PB��H g�$�"f��_�=��,�Q0ދ�n��F_k}('u�\{%���Nl	>cy�rJT�q�(���Șc6p�c���D��r���K���ؒߌ5�N�y��!����0Gd�وm�W�X����uƊ�e��i����;F~V9���&0Yq�|�7Zdw�P���	�q��?+�<�8t���(����/Ϫ����&��w�u�#.�T�a��(�#p���/O�x�����IN��s�qE�&ƪW�TH�Ddٜ����m+ɏ�*�ltԝHl�BR��\��h'7�۳�VF�����x:�ح�2�]�_�޷L��P�����&���A�!�7�Wt'�7��%Rn�nOj�v`|�x��)+�F�dᔶ��Ug��Y��+} �pS�(I(v� �F�^HX'��~��]Hl�Mv'�M<�p�aǾ�����?��.�/���SZe LKM�7�Z�@�����C�=G���0H��>�C��K=m�s�-��g	m�~�n���=��f�!�{ȸ�g�cM���Z�oY�lA������1�r@�t+��/O�N0�(���RD��(�d~��A��v�/�ށ,����w�����j�ktix��t�^�⽛�Y��ò#wXIy�i�����/b�An��d4�s<�WJOL���$�jq�c,�{�C�02W�ႀ��?��3x�u�6;�������ᤩ���k�o"/
�`n�W�� �&09*#S�{{J�;���	i	U��Ne��7�	�>��o��b�Ȭ�x��B�f�����۪���� D� ��I-#|��S�C?�?H��j9EZϥx�2"	9E7?9[R1w��E��t!Eju�d@���У���|��{5g$���gi(^E3����c��@�wnvJ��]����賂J�� iY�A磖 ĭ,=��"3$g��=��n�O�_aV�5�U���j"�k/㡖�v!�8�X��j�Ul�^֬:"����v�)��<��k�����X�Ҁ��H�X�NFg�&Kl�:� yڮ�(a-��Ɉ����y��^���#�>�d��U��r�w?�ާ��Qki��85S	|,1��3���J(�'��ә�^qyU�
���2^a����ϱ��-\��ělh�q�R��HPg��9���%�n��Qhj8��F`�������H��a��Ҷ��un�V�f�X������vH�-���^{2�����}3�]�f���B��:�b�S�`��D��7Ǘ�oب�R�%��R����æ�/G��yr)YW8����>�>�����+�m�:c�<TT�7���7�� X�i*�ǗR���<�+�s���w�^�HR]�L��;�ug&8z3!nNVk+����_Ԏ w�d�Ht!i�����Jd��4�">�K��@ǣ�PnE@�"G������%�����ƴ����D��n(�-x�"5(1�� I��=s�L�QD��)��2�idg	����$�׻�XT^?�a.s')� �&c�51���Ļ�(�@��64�F=r/�Y�[��� �?��V�N,).1Y��PwO�A����`�+W���C��Y�S]��r��;��!@��:';\�~�vѾ)rIPt�F�B�=�.t)�ll�'%qUwU�GӇ!AK8���*w�<%	EEA�,�q&�Jm��^!�%{l1�#��L���6~��6�A����`���9�Q��Jｨ$�A~]J�{M�d�JԡR�h���wxs��"��1t~Bk�c��z3�)�8V���]��-����-�c#zI3���)�mCj}ޥ��g)&���x.5��T%)*��j94��{Eٍ�
j�$�:~�E�埊� �wys.w���bױ�φ���]/�)*O��I9�ڀ�����F�����I��{��E�zm�
H��F>b��јHI��4�"	��M�{�[��t�|	U�t�|�U�D�O�W~츆�FH���`��`xUpR����I�*���/F��j+\�*�\��rr"{m�C��)���%᯿ߌ�|�/��(�J�'J��ȧ�nm���5c˸���E�K���p���SSmOޖs�z�Nz�a��N��P�*�9�ii{z\s)2�~۽/�Ti=e�x����1 U� �q���@[C���Pv�!�7u��)�����*jyDfGl�x�5���x�`�&��A�e�]F��������Y0��.�2�d�W���y�q�U�64�{P�*HH� 4�(��oH9����{�͠J�3�c0��z˛�=�n`�6p��)E�_<<HEv�W�[(gÁ��{���{w~�g���mH��k��.�k�c�A����Bym#���4��Qme��ݚ�%���[��l~�Uy�r�<dP�P�?��k�e��R�nJ�F��1Y �I���芼S�q(�2���Pv�Q�G~�BX�ߥ��/SG#3':���`�_�j�vq�:�n���Y�r���|�����#3.Y���Ͻ5^�0nj�:|Vy�wc@�nR����xO��3z�N�2
�-����ۙ7�T�^e��ᾙ��G-���2v{�	���fKn��bb�u�(�ȩ�SX�u�:k�Ȅ�0iRc�=���)`���aw]GFS4�xS�H_ѸZ�&|G�A�eI�ǰ�P L�N	R�9w�/9G�g89�m�~9V��zrk-?f�	|+��d� MMؔ�n���P�:ey'�J'm�s`Db��u.r�yp��Vm�;\�\��F(ӎ�_X��´� #�6-��$�1�-)$�5���ǘ����qSq��?�:�"�G�jFklD�4�	C�.���2�ZcJkfڧ&ۖ�	O��+=�磟��¬C?Aq>R�����W�H���$w�r��{��j�>c}�=�G`}7����G�_�a\W>���БVk���x7-�,�a���a򦒦+�z�;�_��E�\�{BN��P�p�?�NH�$vK� �W����w�T��A�d9����R����. �(�d%�C�ڮ]:$lB� {
�v��*I�s Ʈ�O���]@6����q6�-ϔ ����Y[���F����D틠$��l	�ӿ���7�!� #�J=p^;��i�j��ZוT��$��Z"	"a�2N�EG�|�+�#e���Y���o��BK�L�p鳻�����[�����+�ǐ�$x�7#�1��ݴ���V���^�� 5�9͒��+0��S��T_�>�'�zü�����E~*!p�:�hE�����E�kmJ��^�(o��
�5��L��(��>%���P�#�ĆH7���Z1����3�mZ�*:h� -P߶z4��,Nm@K�r=ӯ�����ΠM@7��
P<^&p��Ny�����*��3ʓ��q{�ryF?��`��X���A���{Z�vˠ�����ϖ%��׵�s!s�h[�F3pW���%'���z���DC����_Udd�د^8�ʬ�Z������G�+���Y%���z�'�[�J8X�80)�]�����_�[qG��>�2g���}>�\�	�Ii	��Q���X�AF��}��,c���,�_Z B#f�Wj���+Kf�����3i^~������$��`���|c]�5��nm�ȹ*�u"��B�3z5�CAUԘ���(j�d��md0�]�O��b�B��%/���Ţ�!�@�� ����p���ں[`$�߅��_���V�ɼП�k�"Ļd���ǲz����Nג"4��b�U���J^>�����==�@:5��%n�c���6�ַ΋7��^N0���6��F�\fI��ٺ�b�cd�P��Nz���)�E$ߘ�[�~��Ѽ<��m� t*�S��`�[Y�l��ٮ���?FwL�L��m�l������Z��{��}!(����$��P Vf�Q?��٥q
\�fb�����!�
�4y��*���b硊����p��&�_�ks1�_GJ�g�
��-�����DnD����4܄�O��>���b�mW�Y��,�
Mr1�>�n�Q�n���M{	��:��s�:��9M�ۓ�II�1ǃйV��L�D|kW���O�d1�~x�g�gnd���D?)���gְ�WW7��.a��%m�
v*^����t��Z��*H�G��V���`�&��r�;�>�RU�l\��(}F9�OkAwJ��U[OEaԙb�DT�q��cdJN|��%xΈW�4/�H��*���p�\��h2]`�	� �)�M/��ڴ$Ŋ���*�/}@�V�.�iz_>����@�<���Uѷ��qN��1z	\��Ƽ�"^���1S�\����j�Ц8�j2��/�Z�ݲj�;x��7y�������jo�>����f��X(�������N�2�~DG�M�C�%=y�y6C������x�.���C&W���K���"s�i\I��{�?�\龒��j�)+�!#�A����䳋����Y 郕"�%�b�݃p�`[t�۪!��  �'=wJޛ��9�|�F�Do`�;�Mp��d��X�dɕ�����3�`��2����Ϸ�������9؉D��h
}��ϟv�SH�vi�W]qf�>�S�������L��A��"/��7I�0>�3t~��x<�ֽ���Zg��y�܌����w��,�)@�#N.M��/C��@J8�5m�'�r5���~��ih|-��������!޳e��ݿ��;����~f&Kbt��W�B��3�V<�b����܃οV=�e�ڽ�^�:��Svx�]���kO��Ρ��o@�A�龵H�́��0�
Y��7o�-VC�0�#�b��:8级�U�6e�o|�x�f9��I���~�+v�	����!�Y~.`�#<ڄF�xt�&��~���^0�+�.�@��oǱ`��2n�k�a�U�TVw.��'��,�\�D�Ӈ�z{����6~�j(|�;��%�;��-t7���L�$g�Z�>cJR��#��>�?
	14��~�]·��M�����&���Uғ���(#�	Kx~�<��x���\���7j�w^��-v�^+�8�}r�v���8��5~�V�Cq	��
�n)�]J�Ly�%�ܧ���;��'��&�xţp��T�Kc1'+\6���K�}H�6}LL��M�N�TL�aq�Fy��9�40툔���	���!|�718���W:{ȩ��3�AU�L���|v����/�j����O�	� ���e���'��P�ƒ�"5��f0l��m �:�7�N�r�"6ň�)�o 	�yQ�'QZ&B�,oʏ��@�.���#����]��pq���<���ݭM��<%{��]��(3[��bdN�F���$%���f��؏L���3�ܠ��޸̆�F2�q�3O�6,܅9F�����3g�kw�;1�	l��op��	Q_�V��L7�@�ۈ���3�-S��D�!M���mC��6߽:������+��s����F��I�XJ�1)Y�z�����v=^�&�r��'�1�s�e�W-��^}�!&�a?򣎧@�����o�挿���/	��Pm��`^S<�ަA��X�J��~���.�$���߼HY�RߗQ:#`_��SI�O�����g���T�\�3慹b�g^�a��Gw�?����}9�x�2����e�xD\�)#�D0e8 *xM��Y������n���XD�0�r��g�&��@�U8A�d-�����R�)�Ң��B�}G�Ka�����E&Z��t�>��Ϩp+p��]U�.�C1er��O�(�M���0oF��s!g(���/f�d��ߊ�~~�=�1ZG�u������(��qp�k^aj3��K�c�%�?���p�ȁ�\ɬ��T�i�-g�������n��̟އ�}1R���Э������ƮjrGeʺ�4M�ڏ���q����shH5�'PK�w��}����c|ߴ�K�Ȱ�һԜ��$Y�E�y,wFk�
�h�h�Ӭ&�<F}��_-�ܲ�"f�W��#"�r��1�+_�h�e����Nۧ��q�EXF_�3���6W�癒����c�|^�S8����g&Q�x�9w���	�J��!�m��B��Q-!!���8�����r��$1���1�u���KayP-�B:��H�rDFVm���;%G}�X1��܀%�͔���(�ĞP�����8o�OV2A�����oz*�_���JI8�Xj׿:�C2w�����3F���
'
%�&�<�ݻwu��do"�~4�[���Y��x��3 �2�T+c��GV]�k`Z
�ÉA+v����[��9�&KpV=�8	�p�tP��.Jគ�֙���4#`)�!]�?��ϙ��OI��7y�Gn�����`aKl�S�օ����(i�����|2�#7����\��ّ�`�<楒�g��Ui|�����̐2����l�$E^��*k��>@9���-L�ÜNf[��*CS�����������|3PBx�byGZ�����>���Ly����	ü(�4��0`�y�V������H|S�&0�!���f�G��n�gt�E�^�/x��u����:+?�� ���RK�꽖9�4�(wK���ǂ�AâpR�-�w��G�xtGkB�kB��Jo���~�^+��g���d.蟼'���C��*�̯�O&SGa��҄щ�Vi�(&�B��{�j��}*��~vx��П��N�'�]���
e�`<h���)n(��1�<���8_a���݉M>�^2����K�C�S���T�1y.��҈0�7Z�C�p��!|�BU ���vq�� �����e�ƿJY��&���[�JTa��§l�
!?xv�[�ͼ��|����0�b����(Q}>w�оD�!-�4m2�n���Yv�ew%r��"7ή"Gw�B[�hc��{KI�ӭ���5w
|�N�sO�s0����u%�U��H�aj��Ei�"˷���#������6�R�����b-�/��Q�N�O};*2����lCO��U�u�%)��|���gZ����iS6ǣԋ�K��?���k���	q���,u+D�ဋR�Q1�@��3#Ko�:*��Kc�e�
�ϣd�]
h����7���g�1?���������@��w_�)�Y��/m��8�`�4i���l��Xq���B�h%R���7&޽����h�˜�-�F}���k'9̄��3�~��.�j#�N�i�"��Y��C�P�GN���@��y]���Gu��2��%����^奉3H����F�{�avs���Y!*��@�s�mK-�D�	��?K�M��|Zo���f~�'��ٍNY������~V��;�R�#��\�X��c *Wȸ�zN���A<�@���*Ȱ=�dOd���tW��>�楙�F�д���ה�����(4��`���g7��I��2��`�{�7sX Ӛ��U��梹r�^���;
�^����G���D���*x|t)�P��`�t�&�`"�| !U�eiH�a�?�͎E� b�I�)��fq5�{��?��QȐ���MV�B�T�z{ݸ��D�DC�M����M���^��h�����!�;�� qɺD�Uc��	V^�sf����'��{@ �Ѣ�U���]R���)EsM��T�>2�od0E�֫�4���e�1un�A:`"�������+��:�<�/+S��=8�4+�On�p5:��ֿ:΄J��D��� �@� d F⬯�`|l
���vJ����n�.���&,��=��C��a.�ּ>��[��F@�+'��2^�V��1d���u�W�#�Wu]�Ф/2�"���P[b0�^u)�&�P���ׄ*��c�;J���7�W��4��h���1O��0�?�f	L���3�܀ۍe���u�a�ʫB.*�8ϢO�늋׺6��Ia��E#�#z�n���Ԁ���t��D�n�։��	��,w�ȑ���%^�m`��˄ag��ƛ0y�C��
	k8�.~O&mQ���1��
�=p
/,SYF���$�M��y�o�ތĶOc����M݀[>ǰu�c�b��5W��;�����,6�:�0�Y���0n(��]�)�a�gZ�W��������0����0�]DP!���"�j�t�˫��Վ��(� �� ��J2��v�ֻ>�=������,5�����'#��(��llk�n������
�.��������ɵs�5��g�l�F��Zz��)�՞��f�1���T��ƙqťك���w�	����*�������ɪb���C��T�t�X�}m�ee����~�9W=W�X��=W ɧ�t�6v�C��::����$w�����O&(+3W���On�(�`Ω�
a����|���2��M��Pv�4�w�Һ�A65
�S�M���d����<��1�H�W;"3[�R���0�=��Y9�-S9�'S@�0ǘl?A ��Z=W��OV��[7�^O
��������p��xy�$��Jl,���7o��Y&���-VĚœ!+�]�_��?�L0WJ��\f�Vz��6.�\���<�)q�q������K�����-���}FY*>X;��3��J����j��]\5�����u�Lv"��_�W������Rr%Ҵ��gfN�1�sdBR�\ژW$��r�����:vս��r�U1�]W��z���vn5;M$re@oKu�S��p6��^��f�&��{ihz���`Q$��;��.�y��$^]c�GK[y�.�O��7�P�!�	�͟���]�r�����((=cC[������(���+<���|c�WGl���u���!�K�x��!M&`^�����M['1�Q�z?�[dA��!�֖�x�����S��D�$�D� �P�̧��ƃ�p�꾝�L�|7Zay�*$�Eȁ.����f�[��hOo,c�] �ۗ�
�`��|�w�wn|:,�0JJ�λ��`����u��N�Աe�[�5����@�@��]h@¶������]n�B��K"��?iVސ�鵏y�$Xx �B���d����Y�4Л��2PP44$4�S�{�Gp�B��7f:�6�^Hu��D�;9?@Hi x��-�:���w���>��)+�)���'6�J�wL���0�w�?meg��F��֍�����e+�M�KO	��Û��e`�j`m��Ҕ�\�_(C��L:����T���,��t��8���%~2��9�?T��T��T����`Pn�v�?�ky�]@�W�Dǲ�4�m�apqeIJ���#T��H��Y�Z�oi\����q��p����rcf�`�Y&<�?�~_A���㥡�q���mv��
���j�F�x�+���\�i���S��N��~A�y�vƵ���/J�l&�0�R݈&<�k�ogH�NZ�lKQ���Y)�ϖ����R1�<]3B�fH4�*���|]�`V�����B�� hGU�=��槔�	�Z4�9����߻t:|�����ou�(
W�`X���P%�nƝ�G��[G�����RD� 9��#�,��d�٘ߐ�]Q����_�[]�G6���p�
~���o	ݽ���߻=�U�}:�CV�4ZfS��f�<']g��5<]�_��1�~|��߄M-��~�����"��PX���	�7x�����ɠ��ZҢ�@e����R���N�$_~	�o^_�F@����-^�/�v<؀"�j�߫À�XX���N�EĂ&p�R+Ǥ�Jj#%��4�oa�t��������юP�,�s�wO�����}�4�m`���5j�u�T
�˄���O�O����j_���ֈ��g�E��Gm&|$n�+�p�i���`Y]���JO��^	o�3k�%U1�	W�.�"��Ё�x���h� �o���5�X^J1Uײ��U�� $�ݜ%GO����K$��X��:N] ~2͐�]E�%) ����e���	�?.�'�v�n���b�zlZ�Ҩ���؍Y��f�q�iƃ�E�\���^�:��%��ve�#UnAp;�-��t��|8�\z��l�����B���̄>��y ���-	 ~�B�aQ$���>�ٳɦ05�^6�j�<	7Bܟ�0�=���O����}���x�!�B�3[?�c �������2�k���'ϙ֙r�};Ȭ���H�L��tJ���M�J�=����`|ӫB�&��!ln�!�qCm`e3��*X�7���	�ߪ�J}i	��θ�P��C��_��##|5?�OӜ�}QV�/��/��� ��<[a�et����'qt�z<B�y�μ��im�"�I:#f�����Rr��0 ʊ�ǻ�PZ�D���˧�M�e�|��Od��]7U
�Fe&�b� 1G���m�]��-EL�X����YO��E=
'�I�3M������@�=��4A"��Y���<]��IfI���gB�R�1��S��JS���IH��pe�#nLim��"�,j��-�ץC�&��Z��0'�H\!�\�-���ɱ��m�R��Y�;G+�2	6�J��ܬ'�>7rU�e|�F�b�rD,��y V:��f�bⷡ"�3���D N^��P�ZX�������n� ���*��Q:��]��?c��rc�/򰨟A�ׯ�}5Q유hufb���:g����7���`P�|���an�Y����X��砠�%�(����~��'J���I5,�6�E�c�td"�����5T�~��`-�!�p��-m���+�����s� ���m��^�@1W����^VMɽLO�n�zO�x�0�rfTQ���W]�����M��q�	0��-s�D��0�M�gLa'��Xx&}�d�Z��ܟ.`��N!}�+~���n��3�W��g)�]p��P,nFȞ���PZ�����d������b !�� ��:�sC���L]�?��m�٢�' �q��P�ms���T�^��SIK�w�* 19/�U��+_	%�&Qk���u�E���"��e�ˏ=�V;B^��켌PFȏ����dC���z>���'�yJ����Q�(�L�<���D3����.fP�~tv	�].ȴ��uC�2���g���J�)�,	�!,B2������6}���'�V}x��rR�a�z�R�-=�!nwl�]��n���2�"U� 5��K��K�e�|�K���c��PB�-q|S��������P�ɬ9X�� `]���	���Ӿ�W�&�/�$����$�� ����-�zH$I�܄m^�e����y=D��1k�A|��E�.!�9�{�k�+�X�ڛ��|D����a~�����X d��)K_�?h�CE�'��}�8��=6X9G�2�n'���C>�T�~Ӈ<���[� �9F� u_de$Wz���4�L����c���C����&c Awi_�٦������
j�Jg�J42rސ ��$�;�w�zJ,�!Q���^�C�o��L� �0å�-�Cr�w?�	lԒt�V�Q�ųyÁ�9 Γ9�e �mg��Dr�Ԙr��^D:�H,�8��x��K���>�t7(��P�������;�B0+\f���Z��X�8��������:��J�]5�i14��GRhJ��
I�5� �i�����z~V�?�f�L�ۉ�"�(��n��0�����W��������my/$�)��ޝ��0��] �HJ��z뢥�����R|�����X�e��0Ui�_���1�vPw����o�% ;�kO���9l��}m��S����K�Nؽ��q�p=�s��q��Dg����O�}�D�"2�o_�k7�q<-F#�C�c�@f&층8�25{ȿ�os|%��47�X
��/�8s5�AA�QB�b��c��Ik/�o!�����c-��"�q�>f���#$Ep~cq�?�� �j������/��(�qI��ef?����~\5��)��#4��y%�����w1d}A[�N�hy4��0��Hg�Ж����J����"1��s&�P~=�cHl�/�����b��:*��a���H#}��������f��X���n��Eu�Y�N晎5(�P/J��7�M���p_�jם�V6so�NkI>8�p{�س�%�%ju�v3��e�N�@U�)�ɜ-�ϛ�7��1�?s�%�3�@>"�t�o���7n�ES��J>c01�b�\^� -����$.�qXT���C�<5����?EL8�v�T`��=�ąװ뭴�pp=O�]��8��<	��JҤ؞�d�}���~;�q�(wv[!J11���3m��������Z�qu[:B�kI���tO�ި
�D����K$IB�ݚ��E� ��N"xp��a��>U�$v�1��'�1Gc��?��h��*F���rlr��G��_�U��+y��#����azO۰t�h�g^W�+CN^0��}wu��kK"�(�_ce��m�+y5g�)�T(!����L�>�[����I*Gg�%5[K����۟�Y���p�8�Sh>�ABe*r�{���k�%Eq�������E ��V:/F#6�Lڷ��E�e�ԏ;/|,O	]+�,|0�^�t��'����$��$q$m���rx���e���'f5�KD�?�O����Kl>D�H�������q�Gu�6⧜�Ĳ\DaȾ����V5s;cY���Klqi�,\Ǧx�p�/.�p���q_�}�B�p�]�~�8���Ӂ�\]w1Ġ���K�c�= π�"<�6���N��[qMջ��2g�I�iEt8'q�y��%Wć?�>��
��_W/u�HH�j|�
FL6)K�ż �+�aĨT�k�|J3��LB��w�-�5~��[߮fPdC-G�A��*#O'd�G����\b����5���4^�X���<e��J�U#<�ZZ�C}���?ً����� �~�=ȟ	�Q-)I�1��:e��2m/�[Oڵ�q
�Jck�{Y�/x�FSOו��fNI���8m���ځ8`��˭��Q��d�R��`�Tt��t�
q�p�Z�a��CKy�T�L���tZ����d���"�.�A̐�#^~�Q���oV�����Y�)k���C�,g�둃���e�L�'i^M�Na���G4%EP���K|u�AE�3d�z�x'%��QI�:�u8�&K��Î��ky���@[x��'��8o:D�5�n���#��6ܲ*0<�N�!)��Z�3�TA�Hky&��0iʦ��]I��d���b���}��(��#~z�l6�e3�+G�c��{x���o�|�
���\m#J'4�1R%>�p�$�����W"�yu�~"�O�A�k��~�+����Z�����-��*���WdϚqF>+���TZ�uy�����?kBy�|��פ'����=�n���v��l�����>���� ���ȪY��fY8���d4Hp�> Q ��\[��Э*yˑ�M�̆�|����y�]8B�{�ۯ],��s͆�i�7��0����g���p���TB�ϵ�B���D��g��"0�T�Ƌ�P��~<]>�3y�OU�6�� �j�'�Uk'^9�(�/u���\�hcĒ8��#Jm��g-֝�t�E#�θ�������'�f$����8�L��V-�;ku�밉�Ƅc!�``��$�4�l���b>�}�F��d5��:�=�[��UF�����d�IL�6�D��L���A3B98���%��<o6I-X;�0YۼT,�l%:���e���,������������U����)>h���o�s�f'���\����N	�
�4)t��h	�/�d1�ؑ(;5�m��F�f�ߵ���ˏ�x�Mg"�e���7.bcK�ؕ��Z�3���Jj� ^A.v�$�G`�nsK�J �	Ct�]�f�>>��9�^Np�M	4.���}R�qO�T<7Y��OF��X��oQ�[��l����#�+Mk���v?©
���Q(U?4J�'GR&���UKX�.AlOv�e��B� 'DtI��r��B��ݔh�f���$H�/e�+WjJ��BF7m�2�#ϼza;�`�f'B�H�����:���n�Z��|l��x�0|�XN�J�d0����u�%lzt|l���8�^R�~%�r �5��&8�\-�F�Y��&f���36�Ǉ��i��o�5�i�T��C����/�u�[����]�j�==\9�>/�5P�6'm^���X���[�S����ᮝ����*!i��j�[����ᥐX����Dj�k��.���[��D���-2���+�e$�T����Q��jS+�gT0ݰ�%�߾9�\�c�l���9����L6���M�IpM@5��\]�>8�^CF7�q=t�2VD�������ڻ�*�:��ɐ#WB�q�\����X[�y}h�9� t����,�щJwL�N~2�R���>g��PkE (�����s��:�=�\C�cB@A�;2x�8a(�2��)�轭F �$t(�>�_iz��<��Á�D$~��χ��8��h��Z%�dӋ��	��y�w�U�mK��ȝ�������v%j�1�����%M�%��jIx�����䈞A�Mlj���j��z	AS�F��X�C��=$���[��H������P����/����8����ʲU_/��ŝ�6O�٧:ʐ��:����4��0�au���]PT�VZ��G���ќ7�1d�N��m��KI;�`5s���"IX��AntR��z�dh�M�M5��~A_3]�'�t��\�PE���<	]��9X�$���ؘ�����kˋS��� �a��X)8�^ܵ�@�ZL�vԪ��&5K����D�