��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cЌE���M�S�tw�pP�bSخA�A��Z�B�q�a;�\CZ�8�В&Ž'��u�ɉ~��!��5��z��iw5�a@�Q�@m5��<�{�&�*K�Q�f�W�0���x�S���?�1�i�t
<H�X=������ޥ���d���*s2$Ń>Mpe���}]������Ұ'A��X�.�Q.�h�mj^�s3�3��N��+�~>���,'�N2��]�^�z�X�M�n�'w�â	E��ɝ�DԨvl���TNc�D`���w���е(��s���k��\FBT��� ���0Kbx�)�mO�GQ�LV<>�o��5PE��'}󐱉��
��뎊�UG�����H��#z(�ၯ�W,�O��+� ;�l�q��E^cI���� ��L�'9��� "�&K��̴{KX��D��^�<�S͏e%��.-��D�D����ޚ�����a�#�;1i�I��Է[s^�>]9���4|�H�T<G�T6C��������l�����R�4���m(�MQB��mE,�`�M�u�����DG��hdX�Z�Õ�!�0��hĸ��`
��S��6(��#���<g��9�Iy��L���A�c!߇)���|�� � �|��'�ο��@|(�ŮT*&�q~���#��%oI�r���N�X�*��u�>�⿴1���-�MLo@�p�OnF������{ǜK�7.�k�?�&��3�����d|��If�a���'�O����?�aZY?�n)},������(�E�����$8��������L�ZC! 7�ow�.�ܻ�eA��AKU����S��D��䏽���U�:J��gFg!�$���5�^�˹�B�K����G|%8��,���ð��j���TV*"L�p��>>Q� �a�X�=�eZ����h��'�:C�=�	"��ؑV|�F}g�}<.��,�s�wf߯���Lbp���R;�5���~m���j�*��#.��7��a%_�P:
!���&�F�.>�ROn]�����>�i��8=�J���zu��^��&Ȑ�Ĉ��F�ų���P/� <yc�C��I=�N�`=?yoR��|%U���T��$0��+C�D�=3�#��Ŀt�vtYܯ�5[
e q��K�R��ǯ��s�S��\�%�h����e൞��&Փy� o��%>rv�9k��5��6S�3c�]鼢i�r���O�[��U��Fq�W�����&�ZG��D2�A,鱲�j~P`@V���[�Z{�<���B��AyЎ�&�d���������=\�8�h����L��O�������P��m*�A	�TxC%N[�D0�����\fQf�؁��m�o�+��C ޷��}��O;�+٘?S����}z�7���/M�T�@�' Sv޿�1I�?��Y�eby���0KxHT�\;@�D�⠐�C�چ�.g��7��|>��p��iD����f��7黢*`[+��I,t�V	�H/P����RdOc�뜁A��c��&�8������!���/ӊV���_M�\�f��\)63�(96#�V.����c���84B	$�f�R�x�e�����)�~t�qL�q
�;��=^޹z;��P(=���8�g�;��!(L}�Y MI-=҆�	1m�=�5/VM���x@՗��Q��f�i�|eHS�\Ź.����qM�r"Z�h������x$��尵T�����n�5)�e~N���芚K{���8����C��� �/Cь�١�ц�ڊW&x]�&`�4���M�E)>�5 D�Cm[2�7��8� ��Ն}v�<��w�̙_[���2brV4���jS"��=KC,{�>�I	G����*j�N�%)�D��!h.���'S>j3�G��r�A����C�^���\�V���ӖxM�}[��>�B��!A������V:^�t�/��V���z^>CDssҳF��.Z���M]��YS��0���	dH��U���rȓ�ձz��馝�D�|������������u/�\����bIǼy�"�G�7%�R��e�rE-�:���P����2��Sm�qT�UUFC
��l��q6+I	q�}��(�k����@Gm4�X�jo���	�S ���a�4��5uE=�Ͱ 5W����~|�?QOe3���h�dӏ������5Q̎SID� �1�ޏ�Ϳ��o6�m�^ȩj��I��쮖�)����ˮ�F6H���m��V�P�@ɴ���n�BVY�����$X{|�5�pƿ �v`���;��K� �S����P~E��y������8�70c����J&.�+O���� �i�k�o�6�L��N��~�.�%��t�H1V���3�O|9�%wK'"�aѬ-t�:������z��5!��!VR�ԭm�j�蕇�����`~ng�jC�e�E�ڌ�����=a8���E���$���m-�Ya��X��c�(毠x�C�-N�L�����82�	�%�����,;�&t8
X�
f�<��}���$�f���L&O�H�8����80��q��W���V��^SW��0���%n[�h7,;1�M~c�x��ë����"��#۷�(�:*���˾ݽF��gf�7����d�IQ��m�~��IﻬV�3�y�'�D�ѽ�(��%��,�4�^Jѭ��?�%�b�S��2K]�~s@E+4����L��L��N]�;ʪ9��T�1%n?~������a��iR��O�\N��T�G�ɞ�!@ci�:mD���Ќ@V��7p*��Ryx)���͞Ӏh��6[4_�H�DJ�q�Ǎ�*y�h�K}Ff��&�߭��� �����y��m�QC����"����[nA"#��Y���eU�����\:_����v�D6�eQ�	����"�_a��}w��5i(�I��kՓ8*�]�1�9�K���N�)H��ow��*2E'��AP��5]o;g��(��t%Ɛ��
��*u�
tJP�! ����!9�B���QX����x��?���49�v@�%%)�rqS�$�;j�b���<UI��w,��h�a�Ӛ8�W����� >�+�ʎ��2f�u�֦�!+�*nQ�-=uW�� ��Zڞ�;���LV9"��4�@
 ����n�˛�?�k���'�Hgo�e��[��vK�����W�^j9��P�
�W4Nh��MO�7��������hS,@HY�𵇏z����`u��
v�0t%�)�!���A7����}�\�ɇ�E�b��h�X�S̢{�QP�P��D��=ט J0��)7zY%�h�ch�����E¹����,K�i�?JYC��8Mܗ�תNf,!����V�[d���g�N9@����i��#Y�}�شF�I�R�wt�/<�� �|�P�f����s5�#f
�j���?��:��w�,��i+��>W�*���f�?�46��� `M������?���򢞡P�C˾���!#Ǭ�Y!�G9C~|���>�9�M��l�9,�D@����;��v �f}J�J.B�y�����$Ap���dG� �^��=�����s��u��7ˑ\�4]��D�_K��kcȅ�0����VT!k�_��b��ܖ<gT�@�1�E�9��aY_���VW|�%������J��,�����Ѕ�|>j��r��+�����U�n�ZcB�ྺZ�)~�|Z����/ߓ�gDۚg^l)Aq%�"%W���l���@[�ms΅��}[�!ki �?&�l
X�H�0�`��q4WR�^o�4lEx�'N(����k��d���
���d�]#z8y�*Z��XP��"4M�A[�`�[1@p;�sT�l�on����NT��&�x�]D�ά)�寑(�R20E�|r(�����&��>`i�$#T�k�Z�����`y�Neȟ� �a�`���Ŧ?��h4KHh�B�#��f�`��^�Y��g:��RX{P{mn
d���#����K
@�	:��T�LH������$��x�ǈd@X%���4m�Ky�b}�b!�����7S�ss� �?v�jۣ
겔���0`}�W�*��=�r�9���W%��z�7?�cY��#"+��.���}���s��p���i�����F���y�L�f�����j��#�x<W׸�n}W�����X�'3�b)*�v�j��cީm3x�@�HD3�5	L������fՙW���`�� i�GjP&Sz�uu�)h���WB��Q,����f���Q$AA�+ه������,�� M�����<��T� /�TC�+��l$Dcǫ�ϸ���Kg�������i���S������4�4|D<��8�{j؍�Ŷ҅���!���Н�c�{i�D���Bd�(W�0A+h�Tz�2�\q׹�O=&���$3X`���
��F �ui��ϻ�0w�\.���R�����Q�U�L�.,K2E/R��I��8F�ju8��[\ץ-���O���uMr:��,�n���1z^Q_��Qd�\J&Y	@�m�q�u�+��a���I�^�cn>vA�x$���6���&�(�a���9��͂)����h�q�-���� ^m��
8�1uv�n�-��\L*&����iY`&�R�b��r����b;�UHk�"�l��n�a�辜i��eA>[����3p�����
nr����Ќ�~�yIte���'�^|5❌�M �͙�;aj��dߠ��)�T�z0�'�S	rT}/��z՘����=`�<~�]m85�;�Ս��=�!���Ǐ�`��}�ߧ����H��9�/2&% ��٢:���D,Q̙,xTވ�[=�5͙�	�"��)�24��珸�����5B�����j��v��RmB��c":	�l)S��'��4������u	\JBq��7�iq�
�ʡe�1�W���rh*X�4(+����3����}r�D�(}��|�l���K��"k���HJѤ*Z3��^i���ݶ�EA' ���`e�L���=\�!�M7:�4�T"[�L\����t=�� ���zTqI���'�̠3յ��������,�9*�n�6q�ꂚ6l�I�����C�$T�J�^a6Kk�=�{ܪL�|@�3Jvq�L̕�;�u,1�L�x~N�Y��| ��cb���4硥�����j���1$�n�6����X!A����tF��&��S�a�m��+���O޾�2�ƺ[�@'����W�.�j�8l?��Om��ʱ)>����C�n�	�ȑz��#`	��:�G%�0.{ؖ;�0�)����@C�b���z��C'V"���1S��x�J�3Ɛ���֠����J�n��p�T����1�A�Tl���i���p;����r&��e.@U���a������b�_j��c�U?07~p����F�����
�\q�Z;�,IAD�旒C�T.��5z����eb������j����1����[z��!�I%aD�|Aȅ��!�sLA+߷��H�բ0�h0f�Rʳҷ�� �Wu��n;�J���� ��(:v�RGd����gw5�^�UҴ��-"�"=��H/QZ�:�;���s���s�iDn4����[��ԓ�IsF(nb�ȁ�̪�8�Ȯ ���'�
��pd������¼��T��5�uf��>p��E�=[͠����E��jD�uW<4̮�Z=[I� �wЯr����KH*j�H�a���[�'AZ ��Z���ٻ� �UCfX�ۢ���j�X�x��5��U�Ą�������Al�cQj9��Oz��UɅ84# ������U޹Gj�PA%����5y����[�27�e� "��ӛ�*+��+ME�)^��cۙ��)N�5 B5�?��xH��P���`j�a�P����|I�pk��&݂D�0�����D}wPtA�<P���c��$��W��|u�o��&��)uz�/ �i!qK��r/�*Q���`��G^��i���{iziv�AIi�Ʀ��n����D0��(&E�\NoiZm[��``T�N�]Kı���,ɒj�uo��M�ѿt�JW�4�ϕt�נ�Y}�4�_Y�C��5r���9�
�%{��?����g�Q̇�V�3���i.��e��ߚE�~�!���Ɣ6�NoĹ��M�q稨hﺤM'�`�m�ݿH�]Y�zLU�5�����^��k�Adfzʚ<�a���ݗS:\Ź-|2t��u ��N�P��)��J��i�N����{��z��~Y��P��9��	�����m�Q��vd�����`Y~��wO�p`Z�9FwI�'�E� �Ymy -w��ut��oz~���C��I�a�q��6�3j!��� ZB�S�T�im����D`�B�w��6'T[ձ��Mcȹ�*�(+٠6������#��Qj����}��K�a���S`σ2����z�O��Wǲ����'�^�=t�
����YڄKUd}��Q����-Un��KcS��G��Pt�6�WCA�������7D�6�{��C6��Tt�>Z�8r�Xé��z�g��`�?
��7DT�,�D�!{Dd�Y�=��lա,_�Պ��l�M��G1��-�g*ޕ����")�I GfP���kx$v�g7�.�8�U|J��8/��r����՗'w"gb�������Z��E~%��'�/=�b}N#_���YJ�)��%~��X�U�G+���B���������7�(%�輭(	}��"�=Ջ��?P:$�5�wE�Ml	�Ä�
y|I��L�:���Җ��[D �_����iq.�Z*+��[۾���D�o�|�x?U��fE��F��#x�
J��cW����lx�uv��W�z3�[�HC�y@5hb�U�d���2��F,E{w����HhJ��L�*}�m� 7%S���\���E[9�֞ķ��������6[C�(d�*uĀ�}WX�.Ӊ;c YV�I������c�kx�z�ڴGZn2�Y��,װ�"ju;֡C�R>�BB�������:�mVZ�(��A�����]$_:�m���C߳a�5N.�O���'���Yj��fVVZo��Gݓ@�'����}Ԣ7��܆�Ma?���X_ɠMS��sO��XR�.���N"p^���>q���ڼ�W*b�#�k&Tޕ�D��N{b�Ał')�^PgC�7�^�"5�-��p'���?K��-T��*��f��3��à��kTw��Y)�]�U�:mo~���"���O=P������iw
�p��2'���r��<W�󓼭S`�鿟���i�� ��Dm��m�G�����%a�K�Q����=t.]�
�Gw����3V���!��^]o�J>����Y�B���?&������CQ���=<>?��ܴ���%�G����Lͅ��5�ۀ����~9�K�e���,E��*�)`i�R !��׺�l� sv$ �d5 _���I)��7Χ���{�@:L9ԡ�wt]|��Ai��װ�5_�\r㶵��#��ߕ(��N�ߩc,*��W3m��g�*'=���\�;_5G�xt�!C,�������-v^<�^�`��C3g��g&�v�z_��\!a.�u?�?�\ˬ�&z�!	���:�*��8y�;��`��2%�On6{�	o}�f�wS��{>HR�!�B�tuQ@�+�sͲ8�ZEct�����ZV�﵌�Pe��|O٭�i�H�,�z�� "�{��x�w��+'9>+�a8ʡ7��v��D�!�C�,61�tG�a�|L�=$F�|��IJ �^����װ��į�Ʊ���,�N�kbc��'����^���	�l�����]��U;p\��&���������T�0��6�	Ax�U�/h^�`���A��e�3��3��ÿ�>ȿ�V��ߡ|�@g%�E�MI!�dV�y:K��T�8u&�-$[葠�O�駥�� �2´�x����+�IK½2���[�zvw�WY+�~C52Ѐ����d����2��d0W���E>��E ݻ�}���߱�R��!�pH�knOe�9N8���	S��t�� i�0�X�e=�hTO����&sн�r ��Qړ��\"�����|�d�Ǯ�X�%݂
��K�c�f����@�v�@�zm�"�f;�@� ��O�I}��L⽁٤ѼNU�-�ix2v=B������Q����7a�� >�]��ڃ��ST�KD�T�?X�_�(��$�?D�l�v�%���J~ԇ���O�+�`]6��w�����/IZ`��nw���v��%�b��V]��ٕ:)$����m�R}ͷv��@<���Ef�W������GIޝ�xV��� 	!	؝�C�"ylT/x���Õ��R��F�D�~�U�=��$#=�!����R,k��PF+;�O��QέZ�;�0L�ο�e>� 1�'�N��)"���"�E�P��aϡY CR�Ika��(�Z"�����VAq)>���V���Io�� u���V�+����y?�$��Ĳ��O�}���C�*�	8K?���j��=�i��>��2�:&V�����w( ��D{{�1����3 ���p��?#xZ_C�R��i�ځ�W�+��:�]b���5B �t*\X7�F��(�螏}p=r��ܣ�	�&�und�$��<�Ij�`�Կ��O�t�#�L݊��ޥ�6U�y�^�?��7�,��B!3������7/1���X#q3����8R��85%��z�l����xw�Y~7��@Z@.$������"0h��qF�H:aR˧Z�h��U߮)Vf��xf�����7M0�ţxv�^�����2�AVZ��fD���3���d�D�B�ψ2󐪅������c.�S30o��Sdo�Q�=�dd�#���4i�0L�㯵��[k���JG����³
�-��<�)s�ΰ��������sd�&��4o[At�x�O���1-N�(s�i�*��Y�G6|h��W���@߮������s�N�L�S��5k�m���H��$\��X��k�ê�+�x�1��Zų�4,~T�|s�kA�+@Oӽ�iĊ�u��x�<~�c l��H�]��\6+C�h]��\a����Ģ���s����A���"
Hd���BD`��^��o�,ה%�@	���*t�� 58�b$���'�)�o�o���"���ݩ'c��m	��+����k%1�WY1zq�<��h�:��j�#��'0�����)�����T���M��uٶ	���,�\,��sK�ͧU3��ΪL���e՗5��X�$� -��6&���^������#"��[��m�#��Ȩ����Y)�h:�<�u;��3��巧R�J2\H e��u������D�n��h���_�ޖ$�X]�&�$���T��S�b�Ȕg�cr^����V�M�5Y�h;aGd���O�%Ǡ Ry��2/���#��@
A�\���=��9^�����b�m�	��N �V�!�R�K-�g�rP�_��.<��� ���؀s�}� 1@-��K��.��h���g�VP���M��F��$[�����B���$Ա��F�@�+�g���1-�C��@.��́�b�'Z�C_C��������j��"�S�m�g9\�&�j���}�#�� ��$�L�Z���?����S/��C�SS(~�s���	\Æ�g�Y;j�V��pI/�?����u�ѐ>���=�3�Yu�>f9���Qrr^��;K\��{��|ܴ(��v�D��:������^����"=�i�Q���5�:�$8��p3�M&����Ղ
��0��$�t��'2��������F�&���~�0��?���C��*Y�MC���=LD֙���ި��R8����~ ߗ7�r��u;"*�_!�Ԫ��R�+@�m�z���3�J���h���C)�l̺����8^AC��Rz�C�F*3��De�� � �����mzd�l����v�#�K��U@k�һ�0|)�O�E���w� Ի`�q-�D����NOB�=��<5��g
�T��YV�4|��m�[_�ײ��|�u�n�>*P�,��[Y��͢��y��<��b��x���g/ca���i�H�Sʤ,06��ޤQ���E�0&io�D8�E�r8��	�V8��tL��1��[�_nhZ���h'ɾ��tMy��,4hul��g��<{�`p:DD,'�g/�?	��y>"僙Ɨ��c�)-����ciDU�|�&��봒�F�Fa�2U^��=���؛4l1>�q�i�����%���0�������M��h�#���lbK?��%���N�9���T3��7$�Qo�vq�p{ʭϔ����O�;odV��cK"�0��Q���ph4c��k�0�E��(��:�r�9P���i�	ņ�l5>�Pr�2�+�/���;��h��[Q�8����Mڀ�/Jxn	)��@��bfq��V&��0�ܬ+#,�������Z��%i����TK���<Y��H��Sd=��2�Ї�/*����c9��`�WꀔLwN�O�}���-Q����P�R/�7�*�m�^���m�����.8�yl�P�� >W\�q$��?��{�����]��PP�Cfx����$)�2(��JMQ@$��SD�0 S���ר�k�H{��S*i��b���'�|��Z�}ZP�,���$.>O��Kh H#�Q#�}���,Xԟ��8��?��Ǜ5I4�9�7���4^gka#E�j#��l~{m/:pV���{|3���Xfް��En�P��++t�{'l������d���M�S*=�
��-R��P�3Q�8�p�נ$L"�w
+�vٌ�[O�������u"�DW��`D0��G���8AzC��[2��JgT��e��c����v�G��
�Nd+�;�R�wޫ�A@3?\O��ԭLжOKs�k�%��\��q��{jS��0�j� �sF��8�@����h�R�Ȏ�$2V5�oV���"�	��
B����g1Zgdw��(��\^�ӽ����b*�haȡ/�
Z���D㝂�S�N�"�*��H��X�x���������!��;�&>D��|���	:M���Zo�Y�z9�F���0%�Ĺ�h������(
{IΞ&��-�)@��D���`��Y��Q���� FG��!�O�H��E!ǋE���v�a����!7�����5,_Jfv$(�x�[�H��jע6�mڣ��\�
եk�;e"n�ߦn��"���vA5���}�M�����5��δ�ݏ�x>mp�x�)�_a��}EV�.�7Je]w��ĺ��*l�1���h���������z�q�d�R��@5"�B(Ρ�*E�*4vFP7��#�u7��5x)�߽Q���j���
ec�tD��Z1�����םs�JX^?D��{/���:a��欆<ʱ�Hڐ)}��.49F�ҠqH?r9#���ϫ��OG���e���޿-MOM3���6Eu?Am8���Gw��.k�N����ĔE7���?\%�����?��<G'~�_^��GX<m�׵r�#�p��
�#�k���W�<��ԭQ7��E��_�um���y#�� �2���-O�����b%Vx;32Y�U��n�:�E�Q~9iy�zͱde�O���V�����@��^�b&<�L|g	�Rx1) �<)��zr��m
�LQ�T�,bM�B8%Ly��ڼ��c�f�8�u�;*�N�ߩ�τp�Kbd�x�k�S�b�M�%ߒ�L{�/4z���r�֦��dF��'���gP�l�a�\�Z`�Q���Jޫ�U�]ǈ.�JƏg��xo��~.L�߯Q�Ny�OAC���j�f�b��Ŋ0�@��v�(�3�߲�T�Tm
8
)7n.�~�F���Dy�K�'�R⶞5�9�ld�rn0Lje��R`��)OCw�ԧ��n�18��{��-��YX��3	�ρ-�>b�w�8�l��Ê��Z<B�L�0�*�H�^�գ��l�t����}ʆ�7٦�m���i�x6A�}'��ق��V�X6�K��Z� (\��ƛGA�qp)#�� �.��ai�~АӦ��B�2'h\���*�b��$|�꽿C�H���W*��i^~�~M� 6$���L]gjA3ڳ;����{���Q�T�Y���im�[��5�,�>� 5o��u�<�Ķ��?��rI���q#�\�h�ٯ�Y&��p�"1_#�ƫkN�*?��6�9�I--K=����W�gH���^�_z�K� {�m�0���A!;<��H.���h$B��OWd�:��pu7P�f[�b�H�
�Q�]���5�Ҵ��CH\�U��Ї�e]X���R�1jݥv�f�o����=Ȥ���N�t[���+� u��$�%���G����44�Sn��$Z@F z�.�;3A\r�Ed���+c�w��b��ָ�sΟ2i�.�6[��җi�����Ӡr�
1�Z��:1�+�]���7������ �����n>���읃�l�3+!sῙ�>�f���B%�,�I7��1�J��]���r�=��״��e1m*��Z�� �U?��c��h�7��:�~�
SZ��@��ؕ[R�(�����d�;	"�*2�?t#r�\���N���b<��h҆��ě~�D��r��f:4p9eP�xd2�bf7I@���ԒN�x7�¹��'���z��%66�&���@מ�����A�eD��Dw�R)Ӽ&,rvy�e��/�-d��� ~_�����2�jF�������g�;�n!��7��tF�8��=*�Z�ʟV��5b� #)�'z��56m�+��Ap��B��\ʗF��s��-�-D�����!�f.�=EP�c^��p���o�)��Da�A��W��z��.཭��sM�����Ќ��̓���A����S��(po�k� �ZJ#���е�j������}rNw����"N��rR������fl�����QL
SFƦ<A_o���1 O{^�p!�K������V��Ty������r��b8k��v]��YE6PM V����ځ�������(�J�!r]��cW;^Q��K��^�&�3��%_����}�����5S���Դ�r�4�%E��t_�� b��E=Յ�O�Y��Vq57y���e96sM��h�5e��=h=3@�����5�����ϗH������ڤ�cU�ru:ԋ��i�:��?bl>��nBx��5��3gd�� �j�j{��MF���M=�ժ�,@y�٘�&�|�6(Ss����}��Q�Wg��<���pP�k�}�_QS]��)غOHU̓����%�b����g�?DI�t���r����M�����?���z�]��6��'�Ǹ�&��_���;'�х�з>�.dQBŚpFy��?*}- 4����+��b�q�5�Ĳ�A���Dۺ>�޵ԛn���rpT�	�;G��x���ͨIz�~�_�Y��j�mȫ4Æy��P�Nx�����v�f���G�.a�9�KĪx+]��b1���Y;�͡<�����:��PCi��b���������sY0�Ֆ�]C~�OZ�\h)%.���u/̕�ކ�@��|��L���%:
��ܿ׳�)���!٫�%���[������|ҧt���[�kѤo����"^��25��1;��W��2X敻� ���*� �id��P0t�ie���бn!߻��tc��<��u~D�4�_��|?Fm� )�,�8�:ܙhLUϔj��
$��C�St��4�0�Ȓ��U���mZ��bзE�:d��G�����S꺧�o\�<�2^|��pX���nC�g���푌��l�"�	���@!�z� �M#�,��:m(����P�N��t��3n2�����N����>v}z�8>o�5Y����U1��^j��i�v�c�o"U�;K~�\.Y�l�c��5/1��icW�)�ӂj�F`����9̦����P.�G&�ZIw�J*4�,���2ju�j׀��pF!j��k�=�-e�E@��NP�1s��8B�\<*k�:M�e;S��VSh��E�l�
�@6Y���x/h,Jd:H��ϫ��\�ܢ�LA��S��F8��_�ԄW��uD5�v�Z����p�P�B��G#�..¤�f1sب�����-��H��O��(��o>��]"�~��"����9X�-�E��̝�{��Si�)����`z�(�����|���i)�B C�y�E�31>��5��'�0S�vbT�RN�M��dCa
%qGqS�E�I�`��.2�^r��|c"����aI�Ȇ�*���"L����7O��-�+׆�u70 X���$�X���Xt��鵤x�uv#��^ś�����k���� �ǖ|Sҡ߶�r1צ�r�h��f�m7�C�<�ǖL�P�݀�r�#/��^� ��	��}e�h1�𺚜4T^�,��|���	�luИNۢ
�'���J���SFs��@tj�Ċ����Epg����C�z�g�iq�k(E[�rH��zq\1��"���� �'p#O]�A��,�b�%.���%�Ȧ��X�e&5"��a�/��L��o�"C�nxٹ�2�3}�U6u���z^D���m������P1���J���Wz'�{s���ǋo����K�'󪦼aM�����1�,	������v���Mc�r\��`�ÛB�u�HN;���be�����ض`:-$����p���@&�w�:~� 㢁��e�N���g�w\qNoȵ��>���ǿ�<��C�%ɷ}R�a�%8^�y�� E9N�U�9D)�"�r�W�oI����#�J�u'�: V�ҷ�+@H_�8}�:[E���'tK����#��mh4�%3=�m÷y�w�v}�	lE%���3�~�}1}u[�����f��L����^�^Vp\��y��;�ϿAK<�O�~��!�:���J@n��[��d��a�#L\=�1ɵ1o�j����@�g��2P�p�z��y>�DR��X���C�0�޹���U����;C|OkFS*��%X� �u� ;]�T�)Y%��F��h�?޻¾䎃7��7�dQ��;W��A�W�-�]�3�k/��K"�p�{lHY���n�}j��:礹q*q��t�<g�b8L?�I���c{��rx� ����B�ߒ9�Lx�������s����}�K��Y,�`�������}fG�ʨ'J3��!�$P6�$ٲ�ġ���3��t��������(�,����O����O�_L�!7�kU5PagkjS�a�����X�����=xn����el.���f�ԣX��������{v�O�BS������صДK��U\�œ��}��l�D�%����� ƣ�	_㾒��0J��Ѷ�jw�%<�?M��y����V_]�Z|H�=@�M}�nZ]�d�EK��	��:(�#��\���C���8J�I+*1��3zU�Ш���kdy�9+�s�0`�Q�0]-T�O.������^M�ː�
3Z�s|�=��[+>��p�ή���&�q��*2�ԋ:��T+����9b�٤�����ArШN*��0�u��!�#�g1w8�1��>�����A���鿳IL�:&5묏t龓���$�"�8������	�"��0g�m8z2�������)����j�UҸ�s��!�S�ў"e�}<q݂d>}��k��엂���>	��y3�К�EG>���5�SQx�]�R:�z�Ov8X�uL�'��d��%A��ʹ7����D
^e���5S���T���9ܾ����ґ��/�؊�9�?M���y�FՔ�0R�Z��GؤrR#v��Iv��g	M�k�������??5��eR����.kM�H`��@�OɌGˁ��>k^�{ё���)d�
����UeO22\�V�kBl$�(,�yt8���=�+��9����Ы7[o"��D��ˬ�V��&��i)�=�V��96�+�:��Tn{I�yv�A7
���3|_��GG&^�U"�Ln���/i`/V
��)��rr@��yoOѾ�+�Cfj9�֢�o����~X��� >��-o������������
��Β.��p�{�@�`��x�����������'�7�9����g\;��Y*L�"��_1�9�ߛ�ѿEZX�"����M��L��c��US	5	_(*�I�	��o���	����;)��ZX�������MG��C�ti�+M�`�t��d @�9,�&�
���(:��,p0tZ�M	wS4un�ul@�-��������7�$��:���vda�y�q֧�~����hf��rǝW�Dot#�!�gXtQd�%*=sY���~]��k{x�+�b�`b��k�D�_�EH�)���c$���e���?'u�Pߧc��."ɗ��D ����R����G�:��)5'Q�*q��V��,}�u���hY�%k�	ڷ��Ȉ�W;<�w���V\�8�@���O,o\��D~����{'��bQ��@+�Lq�Рc@?R�/�֫�r�z�~�l^4W)�����Fk����a��nh��������ap��a�q����'F��M`ҁ~�{|������c��ߙ+��.�1ʗ�#L}���Ϋ����ZP| %�����h�Ȏ��y��#%�R͒�	9��,�U M;=�Y���~��J�#�I���*j��r�Ac�:��i+�]v���I��#�@n�[�}�l���%`���:�䫗�����;́)2�,�J��D�z��`\�(�CR	�{ƿb<M!P���jx�7��j��D:�V�杽M\[�O��tq_�P��~N����Q/��?�ɞ�h��/B��<Ѣ7#�/�t���7.�r䕝�L�$g��{Q2;`VR�N�5E{|���z����V�?�U�9�F)�P����%�e�0�'����b��1=�lF@Ȟ�	�Z�!=����lK��� �m�>��`�_ooڢU�<��N�Q�q��A+O(��ǀIg"(0�|����<Z�!�]� �d�ň����(YUM��Ֆ�#�W!ѫ	���V�Ϲ�T�̥�0 �%�L��Э�����Z�)N_Ư9�f[��Vя�B���<TJ�۲�##��R��T� #}�ᢩ����;	�pd�#3m(��	��������2��}���O����W�Y���+���(nWYW����)�?��C�� ��ƞ�1
v��w��ŧ�����Ff�)��W�7�����7���Lb���B@�AJѩH02��������[�=��9c-VK}�j鴽���$���}e�����/[�d!�?A��Q�E���☪2���-?���x-�:��3S�+��c�����Z�Ά��!`�U%P����:tx��m��~�RI[�r��ű�y!C_����B8;����u="�M?~�@B'W���E�j���t#vx���rdw�PRb���,�%T�̅�-!�?��f�R� ���E%l�~�(�ͬǡ6Q$69�}�&���(ֱ�K��Y>�w����u�ZA�����#�~?>�[���K8�7�J�W[m�7��|����(9�:��,�ELJ�ph_�y`����V9ʧR[���cZY�v��ؖ�3I��=�w�K$� Q�%޻	r�FJ�T7���Y�X��a��n�VI���p��d5�3�_��:�ѥ�&(y�Zy��6h(�D
R�V{B8�#�Ӯt�xJ��Ĭ݌�m������a-�lé�v�Y�������P�������G�����#U�>4��X���ֶ�K��n�9ީDG��� ߱o�r�u����g��(Wc�Nx���:�W]�Kf�fm�F46q�U5��ncl�t��5X1�[��JR�t(b.KЀ�Wrӗ�h�R/��o1�DXp��`;~B�_�Wa���gr"r������lt���㖵L9 ��5�C,��m�?�9(xxZ���4�*wI��� ]T���n����bgn�~W��j�Ls�7���F�a�Yc>=I����EK$z����,J����8�"���	}�\�p~Ҡ�J>�Yx@X�D�Q�x���m힃������p<�T�P���y�RN�̍�z�����9H"��B,o<%�Z���i�m���ƿ�'������'zf����W��-�H��Q?���y��j^��t,�2�eg���y{���"�d�Ƭ3�Q�^e�,��1Ƅ٩��<�\�]��8�/���Srp�"5��ҝ^�T@����xr�i�����7��#����or�"�Ӂy���-"��&�R,ē���,9l،�#�]��8{� �� Gj�v��tݘԒ �-�zK�*��<ru �׬ 4��V�۳�KOg ����W���5k�Kh#[a��?$�����+{��ke�|Yn�-���`'d0�+���4���I�4j�g�b�F?�C:��['��Ph�~�r!�%6�n�h���|��4/��k\������!Ҿ��F�\9�����T�%W �R#��L&�:���@3[\&<���ӽ�&�R�PNx���~V�HT���V�L8<M�TE3���u�CG9UU|�݋O�
����X=��Eж���c���b���_'����	0�` zCiud�
��`^�Q��i�@(�IՒD��h�&��~��϶�G���q�?6Ƿ􇒟9:�f�^ʈ"�D}��pT+��0S�=uџN%��r�Z��88�t2r�o�e+&�,NuA3.�qn-����9H�ȝa����B����l7��y�*{@�M�\��ʲ�%����V�]0��Q���a)mCT�7�����ib�
L72P��������_��},Z߀�U�n��*�~�Л��.1�KՉ��*j�RD0R�}	��N�'o�oe�(W`S$)ޥ�o򭯓tr��PR%!����
xD�O˯{6Q�qԑ$\�M����<8���o~	׶m�P���6��q�w?ZgG�%�_�b�CB0�+])՞�4t�z_�L�^\k�� C�ѯo�8�j�xE1��P1D����ȝ����'� C`J���*�%�7l��؏�(RBps�'�~3ʷw�%ZK�A��=tl�0@�D����3aY��T['pW�\�Z)�1~y���EM�៨����&i��n�p?��b��^w6c	�:ؤ5ޥt9��F��j��^�>A� ѣLg	�8�
�r�k��Y���P;�=�]��ζ�;�����fDrM�:�q�|ӭ�x9���:�u�X����$F���-�C)�=:��w=DgLr�*�����}F�U�������� �W�K����r�ϋ�D�z����^w�1��]#����F�/k��5�U��NB�`�H. �z�t�ر�pn'�F�a�I(����t�Rf�B�P���	������ܟ,��@DK�^��p)�+b�����jtj-V�5؀8k ����d@�nk���E�s�WD��'���
^O`7��9��x>�M�L�F�G�V��.�̙�9}��0 ���;�y^��a�P}�4į6��1�q=r:���v�9�D�,�ڣ���k*!tg'�B�<�ؾuмv�y1=@lɥ0<mg�7�O��(S��t_�z�g���w�\�譏�/i;���R᷂N{NH�������z>�ܔ_V��lYt*.J�(3;��Ӗ��_ �Oh~�-�_!�V��Og�˨ܙs�^*;��FÂ���R:�*-�/_ΑmE�(rP�)�H��Vy�V�0=���U�}h���A�c�C�{�L��B,�'��N�ɾ�]�7�����\��k���ؾӫ�j ����6Ș�[xåQ��n�9��ˀz�B�AH�{*;ü=AW��u�az�U�q�ʤi$���Y�l�`�����
�<�JM,�Q��#���h����Xqd���txO���	�����ۨ�1�R),�1�a�5�b���,׶Av�u��g���ፘ3k�p}� 9�����S���7ʨm�Ժ���RṶ�~�2-���rp���S��<uQÜ�HM˜4�DF��x�K3��xѡ��"ٰ�$ߋr�����|�WW�8�����A�L�V9Hw���=�A{�KB�� ���J��3쮹G���ol�$��X��V�얖<+���@E�2�@4�{j�]����]o'nP�9pJp��E�g)^�qb&�o~'�U�L?�V\g���,4g�4{Y�Pǣ̙R�(�����w�̨*t�X������y]�&�O��2�p�p�����ڎ���xʫO[�$ݽ-F�Z����4���vS90{��+������[(�6��[�&.�
��86�,l#Yr�Z�
R�%��b����O�{���瓬��Zb�WQ\Yu��]�InF���@�J`8����=A�KX��%V��'�Y���~�Y~D� ]Y}+�)Ñ����yx�K��/�>)��fS�n����]6��泑�`e�{I�)�:D	S�ggK��qZ��Q	 ���픨鄮�R FhM�Z6#�*3"��{)�lq]�K���>��@�A�1��ƔſZ���Ͻ�Q��w&�b0����&��ؖ���$���y��FP�f'QKh���E>�����\�EVٞ�qN����S�Ԏ�[�r1�h�y��8��BS��ӷm�����]{zBz�w��k���f����:�H��9v��],{6$l����c�ٴ��4>ȗe�;y��(�Nk�Ƞ*l��7�O�';� ��V�u��D��u�1ׄf��&v����HOrC�2���� /�Z������u)j�{hȄ4��*;9*m���������P)�΃"J�s'�֕>�<5̴~�����y�}�A��ak&*.���)�����"�|C�.�;�f�L@y���+H/M��2v0�x���q*��������^�m�v��h�$z�ϦT�'���HQY����9��W���Ƕ�����N#8�c�y �R��z�S8Y�;H���
���36��J%-0zv�y�bh�J��D��ޢ����fcUq�f}��A#�bPA���hu��eIHl��Ύ�^1��c;�Q�7(��K9��VK�����c�ˡůH�a�O�����ƗY��i���.~O� �~���8���0<�wz�� �v�����
���C��*�p|Q��-:7�k�����u���E��yΒu�8�HG�%N�+�5_b�@M�G��}"�N�ҿ&a~;�(=��Kn�*~?sR��b1�Hhz��1j9wG�?a~�8�/���د*�c�k_Z���O��P��m4�ϳ"��M�%��b�hb\x�m`�����[$1ug�清WhԶ��g��](� ��������Gz:�sMW������f}������Ìo l���ɶ��t��f��{?m�}
+�ʢ(\�ٶ�f���=���9��c�R������u)%�.�H���"�j��_�h���olg^�:���Q��b���
��/2ƤJ�2���r��G�yl����j��=��呮�
�\�AI̻,��n+���ՏYM��K���#�U*I��}�U�5P_#b��^_M������!x��_hS�ֵJk�T� ��g%R��!�����h�A�U$6����?�ab<��iH��w %���f��+e��q˒h�d��y��3��>�̝=3��Ԃq����PIX$˨kK���O^�_�A�(��ף3߭�.�,1BB59�f��zc��J1Zh�|Eή2��dA��u�R��eC|1#sJ�~j�y}�=�(���S���<���-n�Cy�$�=8���k`��,��S����!�*��}���E!�?|>y�y��+�HBp.�F��&1;0y�i��9�]�@�9�a�����m�',�b`�l'��&<Đ��R��TwnE7�%ur��?�嚦�Jw�@�U3Rމ�|n^�M�=�8Q"�����e�n�ї�@R;e�?<��hR�@�PiV<_Dޣ��Ck)Y��?F�_ja�������&F�kK�:�`�u�L
I*�+�L6��(a_�o��n2����/�bvD�
��Vfǎ��"�aüD�!�;?NJxd��
T�H�Zd��O>#A��{������=������N�i��iʫ�וrP�y��͉����\��E�)��W�0�f a�Wo������aIT�xR��<� ���U
I9њ���`@����LR ��(NHp�zTd���ُY����#�Woqi�5�|�0ȅ�V�K`8-ZM�b�(�_N�a�'���	i��}���r�YP�ph���^��ڏw��)�S�>W���tIbsݎ��c��u\�lh�X	)h���H���~!�XWGUw���&ɔ��+��6�2��%R.�B���P���?׭ٰ|)�II�I�4�?�]��P���כ�Лn�r�8���GO�V;[ r����[�[Ƹn�e�����mݼ\w����A(�Pc�!/�w�Z���5)Ԝ���^^�$pg���~��?�2Jp���)�Ŋ� L�\N.�@�)�%�]&���)�_�v�X��
�n���:h�{J�Mʦ58������l������߱-%3"�=�J�[�L� �h��qo���e��/\�X�?�Te=u� ���p����f��δ���m&����/�n�����)�Z3�GR��0� ..9��LwϯH���4��N:+`}���Q㋬�/�}��������V��u���H��ʡGjLǕ��7�\ \�AN��`�a��׆�V�:�>ܤ�P�	�ϐd���xj��S�/��8_d�K�-C�S�/&��L��P��,��D�}��6GO#f��[�2I�w��/�� ����� ��)O���d��U�(��N��|���ꎬ��'�c���쩜N��S�<_�f������Q� �Vo��,t1m�AtG]k��o���A;��'�i�_�N �kƉ���S�?ǎ	�D�v����Vd$2��o�}�����eQ�R���?ܫZ(X mi��<?	!7�o�Ȫ!�	�K��Aǀ�_PR���HΌ��UV�D�M��CC��M@�XA�ҽ�����YK�x&��U&��:g}X�e9��l� ����y� �.�YQ0�ڳD��ˍ�a�Ȁg��]�ѸT�Z�� �ֳd͹���o��%����}���9���pa.�,�u9?��fc>��j^�Q��8�ֈ��E>&�<��C��<�^#�#\̀���!hR
�6=ꎰE�F��B�Z�Y�0�
��{ ߞ��$v��� �5�L�+�!NݗKe�֣J�E��:�Y���H�/ۼ_�iL�f�,L���⣨�����:��"�#�q���T^c�E�'��꫃j�����vw�e��u,7$^��������1M�4� �5�?y���ɴ�K����$ ����m����>0�ֈ��$5���6��R^_A�扄~(���/�lG�0n�SQp ��L�F�(M����&����^��7�p�,߆��l"e�=�O�����]j k�N)~B���lv˲��f�%��7v�n�O�����Y�V>�I�L��ʪ0���h��fc{!�����$U����� Y��\K5���:>$��/�h������)f%����(R\��Ϩ�Hkk�J,ƺ��,�����J�*�-I�!z�׮dV<��/Ӏ%j2d�(�r�2��l6W�im�p=F���������Պ��f~��9�r�]���s�GJ���8`�:R�<U;�{�{�8>���c��E8�=����q��R�o-R9}�0ɬ���� ����h@h40���Gޥp2�����q��]�fn��^׿Rg���qf���'�hQ���n���S!�cKL�dZ�R�,�p:��#Q�Ռd�L����8L��(A*D�pؼJ+�Z�}��q����}U)�'-�k�.d��uX�)v4�m��
v	��ET��Vr�,�r�W�1r�9�m�j���/D�?�r߮ǐ �uq��ŪR(P��k.�mT���������k$d����_XT���Jލ9_���p�mUAQV�� ���@&�NM�2�K4�r!&����w�!��!2����-�5��e)��/Ƌ��(����t^#8P��*��r���! ��M^��C����x�̶��W�U�i
^��g�L��³
�r��]}��!��z�lqR�K��/�R7���4��q��K�G؍k�b�;l%��A�j��Ռ���/��McCr9�*�`����37{�WU�m�_��K� <��o���Y��8��]D%�N5|F�qw������І�^%scN2=T�����A|��)�BT<�;�!_�ύ��}�S7�����������dzN� "�/m�"V��u'�*kC/��J_+����Pc��3�b�}H�f���v�����~��lu=h�-����<<�b*�C�E��<�ʏ�Ֆ�L����Ϊ�y�e�!80��m��ܣl,�Ą7[GPűT�&R�}�c�ẖ���Tx`�%�.A?�ldr�yK�,O<[Dl�jutW&dm,��_JҚz�8`1˟�[ʲq+Ff�;��h�ϒ�|Q�`5�����2�{����@k��P�]����1(*+gϰ)>H9<����}�h~[�E ��6�d>�B�Y��`�H���-��?�W���_* �_�Z�d�T-�	tHuļ��1!��2�� �W��e���^��԰�Ƌ�U��X2.�>r��)����Τ����"���ETПL7��Ox���P3N���}�uk`\��TDFewYꯨ�[���+C��-�'D_�,�%�$Fؖ2��9l.d��f�Ą����׌�aP�z�<k��9��wJ�t\\9�¶�+�8�Q�dr��5�1l������
���#�A�7�1'|qH�͕�t�
$�CD'Ӷ�hP�2z���9S9�/�t���3�I{�b	��P��&�Ʀ���{W̚Rz:v>��>͵d�K����&��>�F��9�[�&�u�*�W�*QֺT������t~o��#'�Uz������f�"� )1#��8Cj�:�y4�ckÏ��HIV�ޏ:W9�Z�LU(�UK�$�ft�A�������<�����W�R�����0�w ��_�.6I���jd�!��e�������ħ����	�ϋ�����s^�D#���54U;'��0+�x�Cǌ�W;|ibC�/�]��AVA#���,?s���_'�A`��(�vБ�Y���a�(٥��-L8/����r��"�Yk\�
��%sAw���L��?�Y���?��u^���f^��y..��-����2��$�"c߼w����Y��o�{��1�I��o]�Kԫ���=���/���%s��r�#P� ���6�4��B2�{u0Z ɚ@l 	\���X|���|�v�
��xa� �R"s�)Âh���⫃��]�2��Ϡ�"Ѭ�,�2k�Y�ʑ~�c�l�Bh��1c�کU�Z�j�fW��H��xN�D���^�czlI�NE��Խz�\!�D�L�Ugv ���=�ځʧpwo_���2sy�Gхh��ޒ;f��9`�������t�F��obj-�%G��a�F�_�ܘ��b���[kS�r��3[!+tq�v#��pح�Er��jѽ���%Z�]Z6��V%�oM��Ry�I lI�S`D	�JRc��vZ�ZCl�� ��5��˿Z=�	�9�R��yۜb��3�b�?��|�0�(���l�z����g �)��3򱣓�}yq�g���)�u����ߟ�?=SꝔ"%��2ɠ�/�Q`��^A��xj�apج���2�$�[m�8J0��S�I����5�P&Z^΍E�ʖn��pUβ�0e�� &��4gI���˕�VQ�3��ce����C�t-/�͒�BJ�i��9�>	c:4���1Pҫ����j&|˵��=�Y�=��W�3��#`ǜ���+�&�xe�6�S輫�p���FP�d���	ȩ�\�������T>���b�.@ʳW�崶����N����v����"�-�L�I�a�]wN�NhM��CU>S@����	�~%M�|FB�a�"-	]�8"&����z��yI�<r�H�����M�MXV'O0f�¶Lq��vh�D.��sg(_H�LH�#F��E]�.�f�C�VxSQP�T���a�FQa(o���q��7a�#L����SjH{� �u�+��sK���l3_Ӛ@Y���Z7�a��a�r�hBH+��#e���݀z��-�v�h��Sӟ{�1�&`�42�������Ĝ-��{���M�]}��K���$��=ә�o�cAl�S�u}9�5���`!�+X�S��;��ng<��HrVQѽR�y"����Ɛ�����d`Z��.�y�Ԑ�{��}�W?��fV����� S�M��L���>�<����@�3�Nŉ�vxlRo��������C.E������C�0$���h��臘E�`ǰ��{��GD��O7�G�K����$�$���b��ry���mV�2?5���܄��<~��I}�Ep���
���+'v��)��9����O"��%����l��;-�L�N�s?H��yPDkIDs���d:�ԕE�6�a�5D��Ҡ[(v�O��g~SO<갂�}�Z�h��!��\1���
PQ;���3 n�v�)셊��]�7KU�x�s^�-�J��_��mu�?}ޠ���= ��B?�!X�~�de�.��+PE^�������V�$��1�$6v�)��γ�[�b�1�Ө���F$]��ӄ�vN9u��Q�3Lyִ��;c�~>-LYpPYWH��2hBT���l{u��ڰ� 򢑜O��u��m�2��]WL;�%�J�X�!�^alSQ��o�EP�?d��$�h���8�	wV��A^���A)`ޥ�z�-j
���y��Y���C�o��:�Ue�ٷm����]�p�MlZ�&X���T�嶽v��B%ܑ���@ f���Y�,s����z�s��Hx��-�irVX�㷥� O}�����쪸��QN/ef�x�x�ty��a)9F5��U,�������$���yD`��lLcz�q��]섫�����>�_
�O3�Kǒy��0#���ju�M�w�@�tx��v���)���rgx4h���w���ã�Sɯ�����A�4Y�+Tv�����\yW������+˷��LT(�^�tjȹtKW�K�귑�T}a1�9E�����3�m��3P����p�[�q�3ߩ�^�#z��qbO�aJD�m�0MhgU0�Z�w)�K�B�� $Q
5�O�Y߭hط�=T|��|�j�³Ը�!4�v��K�o$�j�!gQ�{R���H&]�rl��T��VA��xM?��1b�9��;ð��5��ڲ����)��
�;�d��_r��������T�>�$;c?���H{���+��q
9b\r��9�Hn�_cCs��4�>�i�H�.I"�m���r�h?���:K��4VY��"DO?mh)�c��+���Ѿ+��f�g�:)��Ө��Z�ǟ�������O������'��.�z0� �=�U��.�y>+�<@V�r��Z�FWʙU?�S�2�	[��H�ˮ�>�;N��/����j+� �����G��[�	���a�q>.��K�f�@����J�r|"(�7�P��7��֏\�/iЖ����5�,:M��nګ�*���;X	
1�����kǝ��Ə��ʤ���:B�*�N8�����q����@ ��_���k1~B�p�t�Eǩu��U��S�^�@݃��y���B�Qg�(��9�c���"?Ǚ��'���d�0����"�G����w�j�en��`����06V����3w���9�d��� %~'ȂMP>*# �+8�Y�96X+����O@�{c�|������d��}K�iE;�5A�
�p�MG�[�|�E-(�=�/n����92���z;����F�1��Ϗ�!r?��@C��ݙԻ�����	��RQ�
G"�����T���xӰ��Q1�jG	\�����'�BLP�S���������M�5�>�Ş{�@���7����P!�ܡ=�(�q��C��4ǎ���ρ'0�ɭND�D�|���<�qJ��w�0�R�.LZi�?�iv����L�&����u#����z��������t	�UE�~e�ꌾ �-��"y�>5��p�a��0�KT��Љ�c/�`^D�)O�'!ണ)q}�H/
�5��Au �����Av�0�P��f��pN+Z�G��Hc�
u��}�柎~c�m�RUJi#�%sb�t���'A�f�}˥L"���BU��Y��j*�88�(K\�c��㢟�|� m����(RuV/�(� �T`�y80��-8��-N�����SEq�흡���U!�*�P` �c�i�*�ux�]�T���9��2�@��U�B�&����ƿ��Ǉ!;~�!�yL|'u�s� ����$�2�B6i�X�ȅC�^9e+��m\8rK�����-U�([�Q����-5��}2���>)�7�}��H7��>\4�c8�JU������jF����5�<��M�F�s��8ک��M�tX�St�}O�H��?Ҕh|*��Ç��a� 7̾�e鐦SU�o#��&�^��$��C�c.�aX��4��8FZMN�Z��gQ4�>�vM"�� C������tx�&��q�3�c�4��9����lPI��+��$����� l���ΌE?{U��%�{��Ǩr\:e�3�)qX�Sİk)��iF ^^�./�V�@2������~)F��v���u��,�a�m��VBmn�tS�|8ML$a��*���/�����<�Lp����S��*ʡ�i��=�d��c���D�0s@i�D�ܚ��z������D�fNP6D8|g�E��un�y3���˽��3YX��iV�#,��SX�J���t�-�� ��96R�M�'ӓ�A*����^�&w���J�$wjj��(T��0	\�U%�Ă��a*-���`�:Be�'$v�Z:���mKy���/ǻ�>�T��h�Dy#����%\���/�L���!q$zU����!-Ꮠ4���'1?�S m1'bz�d���k$Â�@�@I[����n�&]KW��`ex�h��S�n��)� �U5	_d�����T O=�"���
PyWɊC!�4�����uK���Q�XB��r��i��P�o�n�̴n�Hv�&�^g��>h�e&��m�lJؚ�}�#�^��P���<%8f|��׫�9��P�uG߻�M�S��o=B8)�;^�I7����@����q��چ�uV,�tٳS��$o��?L\�n+�P09�G���?�J���U�|Kt �M8�����a�� 9-�9H��6��V��W���SUDD�( 5m�S�%P~��30�.�)rӻ UAB�.�u�URI]+ۆ�.�˨h�KJ�^�� Mp��\��u�˒$���� Dk���!@=qcU% ��΄23���|	l�������[Z���On<0@�4��5�r ��{(��9Q�՛��y.%��K�uC���m�n
F�
'p+p��$7Ҁ�#GQ�xL�:O�(�c�j,�ȦE�a{ ������!X0�î����RCƠ�ME�݈n�l��Xt��q��;��8�ָ�F��8حcW�= 3�.f���ɾ,��PQ7�������F�Jl�X8h�Z<8�#��X'�v�E�7dYuY���,����T�-����Zy>��D���9i�CY�L?0+JE!4*-Ž�5:�5W��Y��W����>��	�)(
��ǻ9��HJYZx�z�K�w%����y�$\圲04j�T����ٕ��@WM-yd�~�u�r�����h?1����{��	�>�4 �<$�+���=���)�Xi�f���5=�B5P�
��QF80��ffuov8���QE/�����L85	^I��i���;|ҍ�.���[�Sۊg�>�*�[�&�rR���pR�W�	&�Υ�aZ'��ݸ3�Z��@��J{�olW�rf˂�\��M�YS����]�O����2�!Q-�R�X��:l���
���s�Q��_�@I�Z�:8�v��r(	v��/��ց<��Z�y=�?�� �֣bZ��쇭���N���O�0O��Rd�([�ľi�͗/Q&�f[�n3�\)��K�$z�Ά�FR^M�@
\�I�_��ܦ�77���IR �2Zv�Q�}p����;�����5�$Y%���c<V���a!����~z����2�c2ǋ�,Wn�!r��O���Ԥ%��MhT�{i z�hK�pb��͹hs�҄�;EUs\]�1�L� �V+��)t��¼�Z�WN�=I
�6]��ܶ)x�0�WQ���j̒H������dt5�~b�#Mi2�c��Iր�QA���%d}Ѭx0t��R��Ay�i^f�It�*Z�	͢�Ԃ���"{�7����6	�6��������(]m�nw!��5m59��Mo����$!�5BX�����2���<�30��!��-�a���Wq��1�k{^37-0��?{���7�L����+6ts�4��-�-�"�h\HT�n �]@�,�9���]=�e�gl�ʪ�Z�4g��x���MuZ$����7�*h�c+k�r���,v%�;�T.����^	r[�H>�Iļ&�s��zgh���3�H��Q`��eWz�LX.�� a�q�ӑ�Se�Ֆ\�,�O��jl�P�^g��a+��5h|���r����Q�����Y�����:�gIV�,�r�b!j �ٛVՂ�3h�Z�uW��	�/�X�g�1�k�E*��t��ȵ��Hh8��O�>nf�	l�ʴ+�>���7��
�9Dxjmr�O��;�tM�'q�2; �1�B ��Ю
��(��ȕ�x99���Lg��a�^+2�p����t��DN|;��\��{�.��M�����t͎�m �c�����	c_&^�݈�F��[��֢���fk'�Tf! ����j���wL�R�Z�1�����/�u,��P�H��/��8\�8��(^Q��A'��6�7A����k�|�R�U(<����M�]�syB�d�n���)|Em,@��x�#B���Jy[ � W�	�7�5WH��d�sݤ�Z�;��=��r�
��,b۫$�9u��*�2�hO{����z�DL�&����v��\�A� �������=�2Q\�8m�bs�܀d�ڶ��<k캥M�$WV�AD�ϗ�L����������x�gr��zcH0�\􅸔�1�����^b��p�����t���q��4�H���R�g��g:�`�©
���Ewh��
;D��xLK_�9��S0�'��or4cJB���P�?;@zةyM����a����\)�:kv?.�2ż)��E�`�)�*[�Т[+Y�1���,'�Y^2��2��E����B�zR]��w㜏�[:L�l�"�ۍ�޽����1g�-�_«��%�	�����CK����7;�p�;��?G|�a;eѺ60�
�.�?�:&������C��XGԤ��(�Xi3+��8�-��S^��*��v��k��{E��$�l��o͙��2�d���4��sT~-tS� =ﺩ�-���u"-�����V
�n��%y�_J`�>e�!t�y��a��� �R���e��zxqF$�c��y�U�� �ً߮�g�F�h��3�)nH�UXw�m��L]>�Ζ�N��kB+�������&��b0v6�~b�
0����3d�)�H������6���)��w�Y�Ly��ԂEG��m��~��x���Ziಳ]U���� �I��D�֯���r�H�h��g���Nnċ�Ċ�+�����22a���t,�	��8�j`��:儶��Nԙv:=n�X�t�OwL�<Y>85^)�_7R?Lh���tk�w�a��Q	����N��!�61b���Ii�5݆�{7��k�G��t��/X�Kɺ�n��l�'
�&#΍�*���>��B�����q
�r�=Q�'Ow�(�LGg�;]x�n�&Bp�����E���_�N�~A���m<��{�(L�}-�
�:M�����m;٧�Z�Sf�n��'��͉s��}g'�8��E5uTv5�����^
�?�oQ�!�ۃ3����m�8����-���]�`�޴��u�Sz��R�ՂU�=	��x�Vβ����i�����ϯ�r�L�(I�qWA�(F ��;��>�㓪�1�\��%�\�ŝv8��e��jZ����� 0�3�>S�~=q?�Ծ+�<��Eo�۫#��4�tu?Rb|�0+$�H֗����f�����8�hIq�-��3��<E��8��l�=cñ�k� �}	���!��>�aK�����Mg�n�@U�E��6����*�w3��0=�teK*e�4��/�Njwӿ��`��H�~_X�P5W�u᤯Dr5±��j+mʕ��������`m�V����`g��ᄍ U�Ż�n����^�D_r��emad�Խu'{+P�I>2c�\~�B��:��
�<�ɴ���=/�E
�"c�܌Z�Q�(��F� h��5x��HLW��xh��	W��ǲ�~��[�*�Q硗���ĊO�����C��K�;���1_��F�� ���xzƀ�>d�,B����$��rh�=�4G:gD����,����Nl�BFp�0hv��ԟ�' ��`��uWzP<���A���),�@9U��4�9o4'�U%Ձ�(6���7��Cυ��䀯�!�7�����=��d!,��tpn����Ӆ��#�������O�:͔�]��m�S�&�"�e�鞐��ر�j]Z�b���8S&�EȬ�y>����l�E��W^C��v���,�N���!+��%�Or6�2�Zϟ���cnb-�M�v��9&{��$d��䵬��F�3nlڍ-h�6� �J┏��DZ���
�>�����
o�B�C�8VW2R	)��Kj��)5cG�Ó��8Y��¢.?�k9.#�T��ŧTИ?�Y�P�t*)�����l�,���e�&�`�z�&S�j�?^H�Q7a��>E��fA&`d�A�uM�������3|.� H��"�K�V��[P�U/*�O�L	���`�S�-�]m'��6�g�'�(��.�, �خ&EGzt��\����o+�P~�aNH.Q�"�������Ѕ��*�AAsA����Ct��^׿�X�Nt��Ĵܩ!h�g�,⫉?�A?�����Fi�W�q:4���JR�-��/+�d�r�c1,Zn��T��t���8߀�<��F�$�S��SAQ͔FOh��Яk��(����֎mqZ�����<[��u��	�-XU��zϯ�}g~����W��On���w:����]Ue�ŜAxε�Ehǔ���a���V8�89O��>Ѵ-�!!����տה=|��cͽN�Q��d�9w�E��_���#V���1�滳�:�;�&�<���s�wt	��AzJ�o���@
XZHx�h���{Y��_j����sd:�he?�J�H�̊���>
�Ju���07	|@.��+~,��:�BV!��TAa�е4 �ME:Ր'IT�U��'S��=nPu�q�2)"��7�����,����A��s#Aq�:���J�z��2Wj����)�J�Hq�,��;Y�w�T
Y��3�%,wLJ�����JC��[5��5��eb ��D�~��0�A�[��k�ӥ���#��<��K�=���j���R[/o_���
�hU[kxs��4�ȸV59��zZu��

H���?ّy��8�=wE⍢K��a�E�������eщ:�1Ͱ�@h�e�����KU@sJ̚8j82Ͳ�?D���g�y�c�T��N*��Zg]��k�_t�'�ҡ��|�Yv?M�`/K��Ϗ)�)�;�p�}�����ț3�;����>�g���'1!C�p��uj���~g���+�cy� ������t�ʝ�(��/&!���`��®��T����?WHB8�S��(��y����.��~D:����-ķ�����(�?}�%�֥#bil��C�X7A� ��+󨈋����l�s����R<췪�*&D����z�|G�5e�<x�4��������h�oA�#�d��v��f�@}^B*�t�#d89�h�Ϯ�G��j����\��+��S�K��U)�����vjH ���m�{@F�U	�;���1&وϫ:M��}ez�^�r�����)8ߋ5e�fHȿn���c��	�Z�.���݁�4|�x��V�D�L M�8�8�S��4>L��~?�,�W!���؇M��Ou�C�ė2A`�h B�9g�4������+F8��kL��x�s��@�vV�
����n7o�>:��{�m��L>����Y!T2����a�<��]�v�zpa����j��r�^n��p�y�j|Fru�I��z�Z��6�y/�I͔���q�nɏ	L��4��@*��Wۡ���V�Գ��jC̦� �Q�*h����V�W���$O�=͹�d��8#<{ �d^�l�ш&�Xl���(�0A������OGSe�p
ÐM��x