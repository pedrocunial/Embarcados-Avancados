��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c��2ݪ/n��g�_��nk�I���h�W��|.Cp�js�ؐ�F(��i�`�Ǯ�M��:x[~B����=��J3���x��3��)�{��6d����Kɜ7A�VZ��� �B�Зn���.�ІEj	�Z*�`���^���T���4����[��O��:�&-i��M���qⵊw�BS����#ב
���10X��8�����i��8�R�/|>�!b��#d@�@�G١PB�
���eF)sK%�����.�#Pv��ת����eU�?�͎;���%��Y��Hh��"I�琟���C����<��n��D��>p+;fL�y6%Jz�.�\$��w���%�I���h�}7	������������҂�}՝��@޶�p�@2O��:��� �;|�ǰ`J|��Q8�b�c%��Wg{��<�K ��n�"3���d_){	�{��7��ۏ"�&௱�1�<QʆTh��ʰ��$!H��f[lթ�����\7p\}x�5�XEju+��Y8x��U�r�׀9��9e?�V�=�J��@�d���1�o�T7�m*�؈��7���	�EZLg�@��}������L��a�7�����9w0�q��Rvui.LޫK�μ��7�3���STb�	OO�A��T�ɱ�98����D^���y���y!E�Q�Kt>Gc��Q� 3��	^"���E���8ڒoR4i�����30�u�l#��ۻ�ށ�J=Qir�5��)QZۄI�� �nr���r�A&-)C�1����u�N�t
LU����R���p���2�N��)�Z���@�%	�k;V�M�#dO����P����/�I�(�/�0�ς�޵�Q���0���i�@`/$�1�H�hN��N-k�pHE��W�6q��D�����d���*�n�.��@�o��M�\��Z�[��X�NZ�z��%��U���Y�n���Q4ζIŀ<ڃ����Յ�O�x�kn�3;� �ks�u[��J$5��Ap���l̍�+�j������9�GT�:H-�Hv�;�)�|Ό.�V�.̷����[TR��jc~X�Tg̚F��o��7Lwu���h.K�̠�);��H�#�{�?ʤ3X
u�Y\�Ƌ%�݊?��'�q��H+M�;���6���ވ��lሌ$����}��Hm;o��gGs�t���A���xt찺 V�XL�����~��L'��A~�<� E��D��ہ�IH��Ȝ~�^'�H�6sM�����Wj�l`\Bu��������O��o�1�2�.gO�E��(M�K��/�]�(6�{W�ck$qCv�8�D'+�T)E���m�.L�<�7>�#\_R�w��{g�^2���-��X�S/�`��f�f�<�uU��f�U��Ծ��b��A��?���7��V� �Br�'����av�����2����),�|����`�tx���P6�)���-�E7�@"	hܻ]����=[���9;{.��t.p�7�V�t�Q+��0�_�z�n71r�#�=?ޱ종$iQN�`s1?�f.Wx��wю���[~tx�-��6�PA�l1DG\�ēw^upB*!7B�c���b���忧��(J����kʨ~��oﬣ�^��R���y��r&kQ[~�uny�M�Dghd���h��#�
թ�΀���ɹ��1�m�L��[FۭY���0bw�Y��A�.��8H�f�]D&Y��F�9	}�G�ngB�JSg3���4{$ GI_|H�����J���Ze�L��	�HK1 dБ�l�"��w_X���G��EϪ.Y�t��Q 2ఒ&p R�-��Y(Э�����F�gUD��D����Hd��x8�J�����:D��f=�Wz���Q[ڨ_�D8��>E({j�Ws�����8���b�!�Z�%��M��N���E�
��O-�Q�;97pT�k��$P���\�,1?�<v�y�ǤR[��;Zu��b`�-���S,���A�i�G;g�_�/����4���%��;ԋ�ćJR/Y;�V����7o���p��`��1�񛮍��~�]�g��I(�܉����E�G��F�+Gbd9�a��&k��cQ�<:�e�X���<	���1���9��#���v$Or{�9l����?Ž�@�?.��	����QyY��D������6i�A���YM�[�����A�v�����K�	��W�`Ր�ê���n~�E��@���cFf�{����vyZ �ZH�`�����zɒ%P�����lxI�e����������N�#F[i�^�oaJ/���mW&��g��R���w�x�y_�g%X�/����Lʤ^�$d��s��� _,,Phރ9EA���0����[Լ�]*svo����'7���fv1!-�a�%ئ���/��ᩤ�F��ed�-���ً
薏��B&b��Ĕ��`��'�}<G2d9�ґ��(�\.�D��G��+�?���.ɷ'� ����P�+#�}�B`{_�9����P�F�?PԲc����D�BΕ��[U�^���i�R�,�〿����tv�<�y�#]
���v�m�|�ǀ����#E�Ӷ�sg�q�@�˥�3.�*�*������>�)6FvI�O0�8�8d\��>���&�'p �<&f���[Lr��2P!� W�w'k��r��ݛ3��=�����J1��	��1��4�
�	��[:��~_�mS�+��:5r�|K��5�$��j��,�1	MA�Վ�o_����J��m�i<�����?j˭qp��G�ʬ<�͒J2Ƶ��5����kD�� x/\�3�rf����=2����i�7�����.���g��I�;�T��K���>Nnt騺-e|{]� ��������b��G�h��Fʠg�	��C����,�eo�yޒ?,�A0,G�%�ͥU'dQ�5���v�kjM���'z�0�cf, жA| �5m��1 �dn���0N��xtni� J]�p#8Bƫy� .�u�a��\�_��3�(��	
������	�zm�+v��ݡ��B!�-�A
�/�xo����;���6#Gu�R .feS�$7��<���������Ph��h�<}ٛ-�j1#�BQ�x�����a��\3�Fv�����_��֫�j
^(B�]G? )"1e�͇m�pp��DV�ɢ�6���.�� ���=$�q>���@m�U��X�@	���/�4�sB�3�r��� ��b����~|-ի^-0��CTA�	�5��O�ߺ��1%��l-f��_�\�_��d�E%�	�+��{�"���>�B�pý`��)�D^�F�pSh�:��+P_��]S�lܸil@�x��m��<�F`]�̺�6��/*ixf�n�t� ��A��I#eU0=��Hwii�ȯ8�G��)���k}(�Ä^�7Hj�W�(��X��t�&��ږ�1��
mQM��0Rދ�<� ^�I
�G�`[�O쬖*��2˰�U��F���A���GH/ƔV>.��z���G-T�`�T�5S��w(b"�F�t��]'������-��D��H���!����n��(>������9�.{���fűP�����%d0ZwT���G�۲ް5�$LЗ�?~H_�@�l�|�S.�N���h��4\���a�F��Y_��8st���9�a�]�}�e9X���LVpT�����)�]zxJ�λ����]E�:0�$��N��{"��h�T,���̪d����Z=�N�%��@��1�<Z��.��	�)k3eh�ɡ������'��|�Oݷ��,��
��=X��Y�z`J����lp���7�EÅ��q��,����ϵ�Uu�Vy���ȁ��]r�	E�������X�[�'�y������^��ū��Q�nA��p��U�py:��${�Kl����o�%�(��dV1�$d��8Q�H��fc1�p�PaҬ���v_R.���2ӆ��L�e���$͸�H��=��! �Y���7�]:m<8��,U��̀�L�I�e�����͗�������󸙒�*�:�x;��5tl�im�VܲXRkA�ٞ
Xre�ǾH�3\nބ�z;�g��K}�Jר�2F.;�,:s<V�&й��Hc��������g��x
��St�����Xpd��f��	"���N3DB֣�\mAҸ� ��^Vn.��+�9���\�]�7����X��,r��Uw��U��_���L���H�nf�,#��&�w��F+� �'`�~L�(K�<3��l/P�)�&��?Ѭ���cq1�Ҹ�'��Ե����X�k�P����YFot��fі*jq�0+��:�u�q�Ә��*��5u���L"z�����+� �T'�`��ߩ"��F ��o�4GyaaxlFF=ӌH8GJbNȥ�aF /A]σ�5�?xa�<�Kq:�W�}�mM ΤE.�E�^����������x�`m����s����:��=w�rSM%���D>�k�c�׃n(nP��������
��[%�����4[�����`��8��]ߑ�I��.9�L���j�	C\�s�������u����Y>I����$�Y����qsKs�&H`���M���D�F}��[���T�rྏE�H�%��z�C�`^A-�7�d���$M�S|�y��u���A��!��h�~�PU5/}�j}S�J��)�.xK=|��lӼ|��z=��P���5}���I�m�W
;߽n�� �i`C
�ܱ4�լ�a�~e^
N�mp��
�A���tM��Oi^�-��J���OX3Ǎ���qM�)u��M�)�),B(4��\�_K���>
[�c�v���<ی���[E8W�>o�������a�*~�Y�0��G���Ct�Bt�������S@AD�4K�� �\s.b�b��Ab?T�e	'Nw��Șt�yY,�oI�V�g��@������	쨵��0*����`�eu:;�]��� �$����c~9��W�*t��{�"6)}j�!I}h��T��?3�}Y�O�N�5����l-��~G��܋�:�5y,���.�-�ۈq^q�i|*żշ���8}���/y���B���O@u���N���m�"�g��?�Cae<ϩ~�er-����H���maS�Pe�c���QM���*w��ٟ'���������hx���M�Х�c�[B�T!��IM�2nH��YC=;�v�^� ���G�����i,��e*7bh|z��<V��1�lc]�c�U:�,�HPUeO�
\N6EmG/��y�<Z,G�COz�m��B�ͤ!��T�1����!G$���WQ���X��%B�3R����&i�+.-���A��Ǯ�}\��zU;���&�^	�?%w۔+��t�S�Tk�Î�ȵ�6�0.�J���a� �jĩ���A�����U�)wE�z�j���L���^�(�ln���7��S�Z)��Yv)	7X�^�W1���>4�l8x=�$QP�$�u��|�ظ��IF���}	�Qϕ�H�a�W��R� g.|7H��P�P��M��	U"�y��af�nN���z�y[>Ǯ�.;��Sn�¦ ���=��t�O�fj[�<�r���l��a�ʄ.�ϩQ�Ick|w?SVP�Z����2��G)�B�>M��g�	�,�l]�Kv�N��<�*߼�Ͽ��^'�V�쭦�9y�|u&!�_�az�"Je�hBT�1 	D!f{JI(т���$�ބ~ۿ�=��]��^�� $�F�v��o��L��(�pP�fM�:�yK��*4G�����^����2�>�p1��5�hg�Ug�x��I�����nWn��H�I�6:ˬ�O:�>;.��B��'qX�(�ͪ��-�xf&~[s������ᑕrz��j�:��ؖ�_�$�Y����6�|�ٛ
pm$YI�aе��Dk��>�w�[�yY�2Qj�6G#�J,yZ���O^�w�uP�lm^�l(F�X_:޿B'��U��%D�J�y���Xi� F|���n`H5�gG����8n\4X����h}.(U9��j��vQV�k�uC<���ǐ��V`��D����7d�6�+���Q��H�h��9�KP�V���M��[�] � *f����̉��|]?�%ȩAu:{9鶚l�s~���o"�G=d����	{��m���wv�Ժ��s�� ��\J�{�rW#@n4�S0�@N�I5����H�˃u.�Z�]�J�ɘX92�}uH�!ȗ���A����VOFG�^�����|۰���V��ζ�Ix�	m&�.�>�re�c�:��m��ŭO��Hהh���JkXlwayT���f��6�z���:GG�q�Kg�1ſ#26��^
.�����u�!���e�3��G�x�zk���	u� W�!�]]���4�ĥ���6�tHɣ����3�^x �#Z�?��#2H�y�`kR��_Bj�n�u|�~������ؕҮC�1�ܒ�hC*n_jZ���P�{�r"�Iڡ%�F�U�H7�V�[���3:���e�ո2H�b��B�`�iXSزvRs$��{�*��%/��ªx�L�0W��4`a��3M-���At7��hw����#��aWO�2d������EL/�q���V��b�(�{�M�9������"�^A}�l��ȭ�Z������r�5� �	<*�3x���r	�}__�.��,(|@?!����N�(YXᔜ���7Y��7-�wa@#��v�n��X��x�*'n�*`�DT�7���N�l#�o�2xlȏ�E�����}n�:?䗏q����<�P.؇DЩd����;D�;�Qm�./�U7*v!,,�{�}�����2�sU�F�(���O6MO��HM����+�Y�z$C��-�?r���(��"\�>�����Fx^��yű�����q����v��Oq���L�R}�`!���p�N�d�a�n���c�U�oY����~վ%e�IX&����o����UX���{,�ш>t2$���ˎo�sp�!��F8���[���)=�i��L���o)�Y���,��L��T����c,qO`���AS���cl(<�<GG��@�*֌�B=Z���IO�/td��H䵧���� m��z	��-�g��?Do)��24�tDcV!�`tO��b�Ɯ]i�a"���O��ț֎-v�(�� �;�(l������t��M���k �m��MCY��s�-�l�<�g%�LV���bDs�&i^�ͪ	U�����Û+����~E��4-�����9/{��2^��Ϙ��><\f�.BS�B�
k5��9I>|�M	��׎�ب����1HB��wr�Oº��(�Sϣ);Ӓ�{ݶ�tސ݌n�]C�v�4|3G'�V�<��%貿�S�w�BI9�ߥ������r�0sd�3�|0._��)����LA�_�˅�u�^uՏ歬�ؑ��LJʹY�z� ��R��5Q$�`c�Jd�䧣7 ��1�ǽ�[+n	�s����ȫ�V
�v�0�/ɑ�է� � C���~��8����&�_�&/��6q�L�DV���tb��I�4v%�M��[P�a�p*g�5�i���Mx�zs�Պ]8��5�L�BT�����
M,bO���RE-��E�Z��:Υpဳy˴���wf	��1�
�L�|v��'�y���'?wf$5���������}�"nQ�"9�/�T��c[�{U���tj~&��#I�gON���{+;���zH�J-��b�?����厡]�6>�"���9��ω��Y%'���u��0�������Х|J����Qs(��c�!�P���LZ�{�M�y���5��ٲ3\5ff�myoٹG�u��`��'���� a9�3����z��;�s�'���1��&��]�)���v�y��m����#�����H�z��t^��=�g7��"�<7�݇طYt�`�c"t�C0�/��\�6���v�K��5J�rp]f�̫�(���m.��-���>�Q@���\�r����^�k�e�\�p���+"��Z&��F�/2&nm{�po+�{,���FJB�A��+�վ��,*ў�c��>��,��!�=�̧��cȔ�H�7����&������/��%�=pR|���Z�a6�+�ܞ{� �V�����Z��Q� 8,C(��������'�`��x�_0�C��+�@��Դ�N�.�T�d=�2�p2�3T9'<�gء�ȶ��e"n!^T�"p�-kUO��zG�V�P�������'��5�R���� n!	>�B�V��%j��(�L��Ra�a}����9�X����<�p�w��B¿�[���q���`N7*}J+�홊k�����P���.��������l�+k���7^~l~t�Qzݯ�����Ǿ��P�(1ܗ��;:�ER��aHƟ%�{Kr�������}��d��6��  Vԥ���Sœj��8��qS���1[�S��7�5�=��P��v%a��\�d����x�@ �"Sl�T�V5��;Q�<���oO�� �i�)R�n�Q�0���qӟ����l�ظ���Ƒ����f�d�����ZΦ�D��|�-ə�� ���K��&a�;~u��ĥ�n!A}�f4yz�����1͸NA~,�nGNWl9)"V^�H��ίCb=7a�4�1��DH1_l0qJ��ʜC��U��4��굁H,���Ħk���X�H�T�7)E*f�r���v��Y�#J�C�����[S'��~��nd.���V#G�Ip��E������^�-.	!O]l�����t�G>1��/u��?�����.V��_�#5P��s�K�?��.㑆�F�B����A�h���}�f�Sa���`��ͥ��6���)�4��,�R_�~,sX����8@�t����y���A��f#=	���(�;��7Y�3�&��hP]aC?�q!����YE�ɖ��l�k�zh�U��KZNi Ӆ����p5����ܸ2I���-��Y�\��=�?���y�$�{�ڮ�&D��s� O	+����;H[�#s�:G��`�k��l��8�=D�=�����W�26��U*,�y�#ϙ[�D*I����>J��4�`R�9s,]6��<�J��������=1�R1T=/>p۴�Q�����"|��*ZFi�g��N��`�ZM"\W_$��_�+��\�i�P�Z�T^��}��{�>#���M��רk��X[Q�a���l���!-E�a��l�??��K�đ�|ޅ*�,��/�YպN��W0���ݫ$�$�f���ΒA���Ywl��ȗmft�Y^��BK�t��}H1�5���\������HK8zyo� U.�Ѥ��o]�5��z�7�y͕W,�4�C%<7�I������#(��������d�&�SP���#�E��oeδFF	��YDƼB�#V�K[��,9�,@��ʭ>��e�㪰�l7��5���D����L����>�׌�dm=2���K��9#@-�z�7���Q�v��@ս��D��'x �"R��[�N�
ꄜ*�v^���3���'�����WQ�;:�[@��M�A]Or�fA#�~�!��)�fq]gF��֧��t��(x�
�
S�M��N��W5O�Ɋ�[3�Z'N�J7/�1j�A�C(y8�0B�AWPG���������e�p����>,$i���uS��X�1������.�N��A�3��z
ꉁ�Er�{$�}w��\��|`�֋"���3v�^�_\sp(���#W�+�Ũ�	)/�'��	q���3�Ȏ�Ӌ\�g.�R�V3��&(�s�LI��;I�7���`�y*a�w�YѷW*|��7���3�:�֖˶{�o�<�c�=��ٱȞ������иd��$���P��?I���vN2ء�r7ׅ>���E&����'�Z��O��ZP�?���%�?瑟��:�@�`>�a�7�=��0�������sO�$
�#�3�P^[�A9���'����;lUMA'9/����t. ���)�7�I�[��okp�g
�`��i.�ƞg��V�S�ǰ�g�,�ʓ1�}-��)8�{9�EU�\v�*��p7��^�:����`V���jL���q��+wڀCG�iBP��qǄ�*�>��'�U,� �=0�8��k��Nqo
h/���w�x�n2e�I�L�j��"5��{ah��ʼW)��jo�Cb'Q��T��w���^#	���h2q~~�(�ƶ72�;��r�悞�w�ᖇ�SF��A��bP�hX`w�M�fd�C�[� �I�M�S/#|�c��(��/��Y��?.�5hF{ #��Y�No�Z�N'���mQ[���/��]\	 W ��4�)�LX����þ߭���_-�����L����3A�ȏ(_����N�4iǌ%�W͋���̓�~�Қ�x���`�\'Ir���
�����g�7�o��}���;1j�F|�̘9���l����W�2��[Ӧa0B��� J>��]�c���?��M����ƣF�ޱ�~����C��^��������m'��窮�R9�7z�[;d5	�9�|��q���~��7�^j�F@)�0�zC��q(�a���E�	�M���>��������s�?O��% E;�(MK���Z'Y�HG�E�i����!ti��&$ �h�`�5R��[cQQ�G�c���
G,Yu��^K���C{Ѣ�ZX!m����mZ���-��G"�-wJ0F�N�>���(�;�2!�
m���g���9�m��%3Dp�P�l�����k}W@�2.�D#s�KYw|
:q4�|��sd�ïj36F�u��x�4��L�@��C�t����I��9ѧ�����f�-W�1O�!^��^�u�������-$)2�����0�m�}tܣ#������b��YC����wQ́��,��T'x�?~c�Z,�����o�&��(|bOG��e`�9,L��J=�B�G��J��z�=v(Z���O)�P�>��=}�Zn���JJ���3�?/m[�ҏ.;���U��Z+��FR3%ѯd�G�tZ�(a �R^�w�f|Sq���;}�뇽��y�)�΀$�;ni���޵ʐ����v�jy�Մ�*B�Z��N��P�9�7���<ps���j���ͯ�ZFT[ckV]N!>�P	
d0��m��*}���vӮ)X�bHÎ{�-)�6u�N�NY\�tn&������g�=�|�Uf����Nw���V�6+�I��oh҈aD�� g�yC������SI�<��Sl?��-���f�ި���_-��C�����VWOl6�j9��`�Y�t!��[B�x#h��^�Px�&S�E7���@<�
�/8�$���z�cK�f������g�N��wC_��-�
��87��0��D�O�>�uo�g�C�\>D@ݢM ������L�.3普U\NNp/)��go�s]R��̰��Bv=����d-� yx{A�msЯ����M�ȤD=��+z�)�9#����ce1���}VTqES�jv��9Ī��R�Ew��c��Z-/�u3)ٯ�Q<��m�zn���z��,��e6ռ `�.X&2H�%g�U@���ޚ�G�� =�0��N��(�[RET-o)��3w4,��sv��d�}�v��������y���߲ya��ف[��#FmS{]$���%�m&$�v-�\����"|��HO��uA@9nPX�t��<��f%t���,�K�>ל�s��lkep��Rf�U��=e��`	;�&�S���Ѻj
��1�T���)��LM`��둥ՙ��;�Bx�%�0�^b����O�������ĺ��H�F�"K�C/̻�"��c]^�9T楡�:B�c�\o_��_8�ض���ŗ��oA��4"�֕;F��z<�!���LRH��F���p�X��L�J$ڗ����Di���b�/�^B�Q�dy"��
o9^��"����@Z���Iye��)r�Tr	�dLJ6���|��m�^�4�P�6�1�N$�b.զ���=���$!J��Zv���]#����R9�; ��W�)Y�Qf@��	���@%b���ː�8���i��-��tΨ�y3"����?��%@�ni��ۈ~�<It��Z��lC��$Eۺ�X��;�XQ.wg��+�A�C����(��wPr���V��O9�-5��!��� d
\���):R"�5˒d����&����i2=��r4��������h�JlA�?T}C#f=���S�V�|V79�I?��Ŗ�g��@�"]�2�rI��֔��P�����Kx�>E������2�6�x�����+e�]!E��Ur:�ƤP�DU� �����̾YZ��=Y�R	�.��R�4��H�x�}A���`�>�3�C
ʏ�4<��	���l�ˍ�g}T�=lf�`�
��,&�t��E�"8U�1� ��xu/�п�xi���j�a�����-�O��P��U~0+2���LJN	o�7�8d��\7|�0��0p���1`�j!c���� m�)M�����6��s�z8!��xlA��D����D�]Jm�~,�_?d�1Vu����\�I��\f"�����y�N���z��؁Ŭ�q#j��ɀK��y7?��`�M�oJ�pK�M�H �5�S�a�/I�L���	ѶFj���k ߙ���g�hp��X��Z�J�ĭ(b��Pě7.��av� �&}^9��(�P(�eG����]W��(�A�UBp��*��H�*�mIT�M(�}:��b;�on+�M��!+6ܼeiz���`%��LaCO�o�W����g�����~]@�����u?��.d�&j�UܽY��)����?.���aGT����>^��#���p�]M�[7��Y�ܹ��2�s_}����I�?p~�&X�P���KC���RY�y���F5��4=>��t�Bw"��-�%D��Q{���������a�����cW���C���-���T��N��Qv�V��c?�����M�x�@Ԙ'�&�4���-�GmqA� tE�S'��L=o��*����I�y��ܷo��9�k�|X��jh��}����P�`z����g On��>X*���*#�n�*HZQ�f^O���b���*��ejԭ�pd|1����	��)+�w��G�gh� GPh�J��,�L+8��`@/�z1XOj�˺Q��e�3?�����U�pp�X�����(}�@�-�<JReH0��C��2��q�B��Az�&�}1]#�[l~��i�	�pQ���IHl;��=���\��jr0��4�OV��Y��g(�+01]n�Y����YV��a7��\f���#bj���̍ܒ+�����qpg-�R���
tچ�(���Ug��L7��m�7r�*
�gP�a������xW	(����r���S��db\��W���;����?l�7��v���ޑ�f��Ny�nc�,R��rH\f{�T6Y�[A��NI ��T���N��
�Lɇ��L�ղw�<c¢���Q6\���>�l��K���,^ۄFs�/L�L}����=_��<a��S��R�D��4��Ϡ�#�Y�����ì)�J�������K��Z��%������]�;�g9���T���@�4�ğ�^�u�}v�a8Ț#��c��.�M���D���ڬ�&C�t�mj���E`����vc����\1D�V�#͢�ύd!A��^���#�3�ι�X4���w9]���5K�yߜ�,�)+i��*�m�����ƨ�R^��)�(t��0�r�a �26�5s���u'6Gb2���Y0��i�����'�3A�]^��`|������d���Z/�M0B��d��C1B��V��]��%��䷡�<��:�Yw�`�}�o<�AI�P*^�X �U����.��풐y�@�F�*�����ٕOMRn*�f�/?���F��r�&�v4}��e��L�|�� p�g"�\�(�G�CrNkw1]�+��ao���W_�
$�@�WI!ٜ]D&bܶz���/�I;jȍ���8�o+�U<�
�vT�](��V�_���;��F�rK���&�}������#�]�cH�Q�e���Cu�Lf,g<�*ܼӰZH�
��Ì���
}���L@`���ǋ��������l��$^���w�U��a<�V���O�pC�5po�,-�1�r��ֵA9<�Ǯ�,s>���P��}�4@��d'���V[�}�f��*�WQZmՂ.3ܕ����3�Ai������vH�D��q7ìq��2(�]��Ssy(��2c���_�/�Y�礻!�E��F���)'�JDΎ��4\�-�rt_�Nx�K���6�= �V�w�ր�1F�
��6d�*��&���z��ܡb��G5.����\�ҕ�<̹<L(���ݯL~˞\}��L�0�2���9�p9�������I��HH�ѵ4�ќG�v�y�I�(Vxj�NJ<����@���9��g2r�"!�#�����7��qQ�_�1���-���~`��`�2%]�P����/H�Dqg���Ε�	Q�l����9�5_v!�:eaL�r���j�P���m���j2o������)�Ϸm�y���qvmN>w �&����v-�ϑ��&7����g���gn%Q�nL��R��'1Ԉ���zy�����և��O�>�aІ� �N�l��V�y �
Z ����pVֲ	�%Ε��$�lA�\�3�m�a7����TXt46�G���)�'j�@��P�{�8�,��	%![wl��>.#z�"���=�*ؽ�6���hN;��u�k�>�St���+��ߟ�I7�M*�nɖ�]D�M��G-:gK9�!�k��7Q�(���m�e�U�N�X���O	D���{<����~���x�i����ГR�f`�O�%]�����F��L���!�Pi�H�Y�	>��~�-fO�4"�n5p,��`��gO����S�n�����X������Oo-W���)+��sc�ROj�k?J���#��V��{�a����b~G��i"�����_��\*�d
E>�nV�?嚶���H�x6`�}��H��B�D����m��_N��z��[����
��;�n�J�ԓ��E��v���(U��˗h�0̧�C��;t_�bBUV[B0) P��C������ş���ikNē�~%�.W�Wq'��s�����=ȱ�q�kN\�{��V��'���j���v�/R.�n'?���� �/��4DNV��ɃN��07��Q��"*]��%�&6�O\�GߊܟqxN�q�|�R� b���;��h���O�}�����~��g���Ĵ'4~u 篌އ�LdB8t��l��]�/FXFP�cq��.�S'V��|�Z�8k3y?`� ��'C��0�2�@���5�	�9E��3u��5���ʑ�j�r�l®���2OC�8�ˈ43|���w+wK�u��5@�k'"̔#Me���)d[Ol@a���2�ӳ�󷭖_�x��}��ORT�<]���]*�ӹ��ǦT9��ߧD��,�N���C�*΀��UX9�	f�1�fs��ݴn���X�e�B�~52�[(�u3�L�,A�iO�5�l�<�P:B\�>�U������^"t������� �d��-��f����{Xϒ��`O�l�������z���I��c%,�r)W���Fc�����`@q���0()L��.���`8�>v.x�W.8���n:e#�Q�Z�t�Z6#��\����!˕x�p��
��_gz����*;Ў�E�Đz��P�a�=��5�%�W�(��>�f�� �w���T��	L%U	4	oڶ��j~�)�@�S
�ƽ�"7�98�;��(��gV:�+��|�g[�_(�*Cbg��{@����V�C�H��lE�b��]"<tBΠ/j/8vo���q����_�08�#>т����?~spF8X�^ &�i(�Г�R��3g���Z����"��[D�v�����%_=3f��Ϟ��f1b�G��uGX�;�8���y��O�jYְbY����^!Ӄ��Z]���o��R(�QB2���W����/�p�ɖ��"���ZȬU;���[�뇵��p\�2�I7�<+�����*��� 9�k>L�@^��NzG�2�'���!�z��d�S�s��r �	Esv��\�̊��0����^�*��Ƌu�۶;議}).ԝ#讂#�'��%�J.e!�?��y��Ȗ��A��t���cZc��uL�;u
�*���@t��)[��}�C�]���t�����a�p����k��8P�sd[C9�*��񏃐�S��R��V�����öF����˅C��[|Q�g$��fb#� U���p��rm���}��z����E��6��H�Yb�@��6 rσ�����i^���~��¿^ޤ��9W�Ԓ�M]���E�6�]�a~�U|�z��'�Hgy��R�	q�*�3�^T��T�h#[�^��� ���6�Z�@ZF}�9s�C7h�$��uhT�-�#L8:С	��yQvM��!�Xe�ن��oeGI�����&1���X<����?9AbCͫ�Z5��!����RĞ�����)/�N�}�/28�F=�;r��ӏ=3x�w�WO���&�.�}�������+��2���mB#��'X0�/��G�%ߦÑz1�G��֭�?�=J^S	e,Ѩ����V��"�kx�~,hP��ߋ]"L����-H�9�=s־�����T�Wp|��H)��}��%|�
J����@j���Q�v��=�	���eW�Z Y��M���ZLW�
�ٟr-����0�J�b�l��c�M?�	L�k	���U����
lP�SX���K�L}�Ț"��?��I�ۉ�KL�-K����.7����c c��[�J�5	va�N��,�Y/��Jf!_X�d5��{Mt��b5���KAx�)�$�|sZ)�X.u����Xҩ�}F�������*E!R$ʄ�V{��i�����ߑ0��ȧ҃���P�)���c��R%k"|6��$`.�%g@�t��DQ�-Z��k~��=�n��� �\'[ݲ���>�CE�γ9����5�~�Z�O�_ �Wݕ����e ��w28������x9����|g2�1��G�(��7oH,��ZLn	��}zz����1G�*�ǿ�7s��^\�X��<�NӃ��ٜ�Z�՛;�w.P��d�W�C_K��Ы���%6]E͇ {R����/a��jɘ2�^�[Rg�M��w��t�X;Y��v��0e֬���1�\���K��raJ�b�@��2�AN��Z�6�w���pW4Ϧ˱�r��k�pM�8�!���!U���<�m;����6r�:�S�z���r8:�Ѯ��Y,X�!T}}
��;���݆ �q�c��գb��E1��P���Uޤq�K��0����g'���8�q�z�4�r��upY�iX�2���锰����xf�5�,3���ޔ$#/�#Kʍ�{"7�G��C�ҿ���&Y��^�IC��0�Ճ�����<����p���[��ƪ��U��5YJS��T"0��g�O���Tn]�:Z.HNmE^:)I��d���9s�Q5�"(��T`�e�l�i���Zz	�!+�-U���<�UE��ང���Ac�X���S��!O��Ԕ)����+H�̾�P_�d���gJG����@���u�8��  �-c�,F��)\4�:��8u�(Z,O��اV��G��2�D���fHG�M�(p�p��$�l2�x7T݌yF\J�ATӔ��<���]CJ�؏�r�=y]�
֕
�G3�ך�ZQ{�����%?�K�b]b��-o^(!qZ���"bY����b�;/E� �U�s���ER (�WF.�_>x��(y���ŉ�HXŬѦ4���k0��h���L�k��L�+�M	T�	G!�Ɩ�Wk�)TM�=�F�(��u]�a���rDb<�O&feX�.��,��=N��F3�/̾��Tg������0�kR&��/�.&�ꛦ`��a��.$����5��������.4Z,�V����aQr�[���mͱ���fJ�a��I~�TOn'��h.��B�A�BCW��ʔ�-�/����7�+S�&@_� ��"����ۭO��L:�-��L��β�
g��D����>�da �A87��Eme��j���,I���D2�mnB���`�C�<-7�o�a��R��	"����/�a6�>��f:�Oۼ��OO(m�M�W�ii��Ϋ.�&�X���-cyz;�r@��R���Gb!.�Lt=1u�B��ʩ�'�Pn� ܏2�J�GZ�)���<	�牠F�ҎB(��]��6�ի2��2v�Ϋ���kSKu�����og�e��:z:)�cf���%%���xkɂ5�x[-&�dV�H.�@(0��5���p+�>pz�����#I#���j�*�F�����)|��>se8��T��9�2W	*��)k�K�	��ȓO�T�*�c�Vt�}���U\��u4�P$H��2�5/�(mՃ��Z;����!u�*��M�V.�z-��(���]3��2!pQ�|�W��p�W��C��#�u���X�{���p�#$��;�h�9���e$�SN�tOm� Ue��zfL����#�Ex?C��4U,����V/�.��Q�(t�����=a�G��#�n>����I#�ӯ�m���d�e�AȘ�×�]:��ʝW�ٕ�M^:�m.�H����#�$�`�rzsJ'{$�O���ד�1&�gY�骒�/��WZ�)n���%�"֏��f���զ����`��e1k5�7ğ��JOQ���QJ�V��U�[�=��r�.
��E�K��ՙE��i�-����}]�qz~5��IU�3_W�[��g��<}�����U�j<Z����
�`����* Ll��B	��������b�����x��.�����Q��:�iw�4ū����Z�P��M��n�����5f]�#�.��l\�>���nI�1�:F��لi˻H����izP�Q�z?��V�KT$�}"�\0Ev���
�Y�)l�zG�Ű���[��\ϭք��s���;�7�\7p���4��p'�!�C-/Yb�!%�z��K�@$�y��7ֵ�ū�j�ʑrO(�����.ߞ+ݹM�Gz' �^t�2�{�]�2��!@PO\cE�ق�U�r|���>4�ql��M�v�Q��J\`T�!��v=�-8�1-yXS#�x!� ��W#g���tk�J��3S�r�����$x��0M����s�@���Vٝ���D���+�`(G��	}|A��~��g�`A!./:��.������ĕBG���?.����D^51)l�IQW��#s"�Xdb��ゐ���U�~���*������Ջj��`n�<��e|��z2;L�Jb|ZCε�0�����[�A9s�V���ct�C-�?[*�-j
D4i�(Ec��ǋ��j���Y�"X+i2�_%�����-%j�ν�8g�3K�U�0��2T��aK�ֿ���8�l�͑{0�t�i�4,J�>8քL?���q�Ys�~�ۡ��&�h ��]+\K�yeT<@����ӥ�c���� {���v�q(?�W�@�q��.^��
�
�	/�WV�G䪔D�9x4���-���:���`�~���ɤ���9%!9.��y���Y�6�>���;��Vt���Mb��t�pV�_�d��4�J�,�:EG�#(aTo�?)*;�M��	�O3��Ԯ�_����EoU��e��lG��"�1Wp֞�!"B�D�Q�b��1��#�!�.f�_N��ߒXHE�1���
�b� �l�[C�wg����7[��J*G�L	X�i�N����r��Q��:�W{/;�Iq�_k|<�t8ޢ��7��[�DPo�+<��I�l.�~}�t�ן���H�Zx+���~��VDN�2s$�7�+F
&�l] +����*6�6ZD�A���&U�*h���e�6��bM�%��"R#�=�`�@EF	���T�ːu�:������6��=�H/��7Í��cm�(��o!���rC�˻��^3���V���-r�þ,���ݽ���uC��s-H���_��f�?x���,�;�uΙ:I�5�s�CЭ�Q���E��[��2g�lI�E%�$pM�H~D� 2�*J��M���_DR��N1��*�҆�c>t=�c1����-�a	D2E9�a�x 薙�㸈\	,����mG���MN�:���
-�n��\(.��g,��<K�vv���fm��M%�������Tc�Lqvp�1� ;lK�
�S�����D��O/���<ozy��#c���[��`ݑ2j�e�j�{�m5��W2���P_����5m����T�u���������Ec������C��$�?�f��ɸt���W���Y��(�}�y�U �H��jƳ0j5�9�9Y�G�B�S�lz��ʻ��_�\*m��VH�."��n��R�t!sUK|M��09,�Eta4����t�ga~ ��o8�
x4������P�=��	��)��%b�#>��jn~�؎'�r%��d�5�cK<�ꡈ,��w�?D�7Vv�y��!�38|s:_�5m��\}�#L=�-پ(�}T��[��j��#n�,��!~m��~��ܕ���2�P���X���N�;ȵ��2���:r-���i�j�v��7�c���{C�Y�@���q�y�����ȉԖp��|�x��%�N������}͗���k��x癧֡��z��#�O��O��vP�� ��ᡔ`�	�3�l߱�0�Y�F�׺�L�n��Rg�Ҁ�j�?2���<b�תn��_x}F@�%oX�F���*/��Y&��yu`E�-j�М�r���XY
&�g���A�odg]��]!�Qu�_x�rW{�Hʴ�;Q5�Y	�I�;Tr(i{�e$z����	*�5��W�k�ʶ�����{q|����|���A즈û�k�7���@��+�W�����%����'�\�[Mm�d�����t����"��7�����*�y������t/�%e�����r��'LUS��"�j{�p�ت(wk���C�c�	�Z�2����2�4��HG�Q����x��,n����6h;E�CW�Bj`߭�16��u[X��r$�z)6'��2ׇ-*�sE��tb�N���B@��l��i�Cg}Ғ󬨅Dc6αh��r߉�6)D!*���yyH�.z��0��ؚ�>�O_h�+����==��7������@m���Lֲ��b�/OD7M�5hAȈ��ac�]�?烇p+)k�~|�_iNb������T$�C�H������`�ߙ����ߍ��Xv�I�������J��fn���{,�R�5�W���2���!9��K���PY�U����FEv��-� �{B锑�fY�}�ޝ��Z���.--��;�*��0��؂�@�*[eB_���/���c�ʪ�G�_�B&���^��e�l'��I��5��Wy1����6H_���l��nX�(��g3��8�� Д߰�ɚ����qEJ�n��-)��ؖN#=������]t�V�L ��L�ېb�:CE<χ��j���"��Kg��v�����X�K�x{0���l^�6��yN��e���[�K"[E���vGD\|n ���>Ε�|7Z��*f2�/u�z0��A
��&�l���=�=r�~Aw��c�~�+�!bu�dʎ��9�z$Qk���u�&IrL`���?��r]U}ҫ S%ш���$n ���8笑�f3���E���eW�f�(L_�y��53���11�8��έX�/4��������~3e#C���7a߻QJu���BE��p�S�Dշ}�&6]`�aBE�T�'�uu4�b�ƧP�Z)��'���"�?�|	�m������c�PB=���o��]����wz����6{v��^i'ߥ�����꺯��Ϝ����W��bnb�r��Elv^��i��rw5:�i���hi��i�tiu�6~xE����֢Hp �O�����4A.����l��%	��W�(B�L5��L%��Q	������?\�"����Ǩ?�����z�̱�9T?Z �=���d$vM<=�����:���5)o�|�ǐL/̈́Gր�`v�	Y�&\?m�"�]���,qb-W���Q�b]�5�A!M���8h�*\�v~�puI5�Y���!W�S]�PR����G�����)z\�����ƺ�\�D�e���7}�="�ā�g�5�x ����X$��͘�ÂDu���-�&g��M��ٗ�Ԫ�A�q�4t=^����#�9Q^+Z���	���\*�}�,�l��:�C�Aw��/^�_o�2��9�}9��m�k봜�+Y��,j������Ì�(Q�p�YJ%!����N� ��n��&܍��bV��L�L�EE��[Zfo�-����ؽ�t�y�ı���ٶ|�0���N ��~�'8#P#~��Π戋�̵���l]��M���1��6cC�K�����Ep�\oj����9���ϕ�a!@V�&�Lח�0�"�'��D̯Z19 D�
�y1�H~�pu!y�N����f�5�����/�E=3�l�HG24	㷋�Պ�>���1-��;�7�x%q��N	�7�����Kp�,ޱvBSLA���5l<?�V�p7��B|4����igp�d�����c��Ξ���"c[�֘��nj��0R3���+�o��k���笆q]r��#�e|n���M}�]=.U�]���טD�9F7�1RŸ���c�� w���F����w�)���+�7wh]6zpo��1�rk�T���,/E�^Uv /���c{��D�˰��&+J����� �Wu�txG�\M��{����UJ���+~|�i���ī-/��@c3�����E��
��-���E�G�i0C��� ��uT
LBE�Й,�%&d%mL�}�����F�zE���͌Q9ߐ��/��ah;"�2�?�_(�o���\^،d��v��0ռ���S͙�ޏ}z����F�3*gT�6���}�^����$^�rAU�4M>��,Ul^�oץ�\��[�}��N���|��.|4o�h�7�[׫4�I�68;M��6�1^߆]�H�-}~�uI���$������6*n����]����v�^݁#��Q*��ns���̋0��S�~�z^��=ٰ�w��v�`�*�Uh%r n�����z� !YC�~cu�#]�DC�G^	��� �F�H��bu
f_Ԙ�&>ag��b��c�KĞ賤��JǗ\*�Fj�ҏ];S{񆛾�⠂f8�8K}�'x\\�w�:�򏦀4!2������k��ᣑy�i��xw��%*�W���!ߛ�����d�XG�����m�>��3������������*�.�Bԋ�	�n,@@͵��4���D�.�<ظS�D	�<&��6{�ok��^�s9�L6�x��s��W�I�J)�t���y�h\c�匤���K�w��+ۏ~�<��%������{����c��B{4LO٦C�E����n-?�[�V���cЬ��|�������@��0|��#���<��,���Ds�#&�����ĥ8�Cq�ݛ�O��L]��*1�������(<�ai���[��e$�HL���z}���w�Joeyʑx�	��%Y
{�;`(N��V��S�����C6B\j�^�7OR�ny�9�7����C'+T��sZ��l��u�J%�W�t�,<�D-|�4 Oވ�@�":�"�)tѿ3'!x@����\����OC(�&�i�X�?��]A�,�k�'N�s��B,PY}#Erp"MG�6�w�K~���[�u��@�rFX�M_(�q�'ë�j�R]g���;����y`����N�3	4����K��C�twp#���|�e�ۺ��>T׊�q�F�����AWB*�1"=<��( ��i�k��!�@48��r��1��"_�H'�qp�yd�P��W��ӐU�W$��8γ��alt�?�]1������,�u#߉�|��V��j)�` �;8��z<��"�T�v��M�^�Q�[�����U��u/�f�"�C�ݏɲ�,n7��Q>@vT��TO��|p캧�.�HKk��%~��!r���P���ת�.��'��Xl����u��p�I7O�tv�G�Ì���Y�޷-�����q�y�.��^陚�q�6$e�f؟����[�ye��e9��1޿�'�����Y��"� �2�?�=T�v���>���������p��E��2�89��4�:���.Is��"���x�. ]�tګ�R�:�N�`b�H���Dg���<4/ф�kO�ZD�$�U�P�{�9>���L��V��R?��3i��й��ﳅ����P�$a�*_H@$�Q����E�.7`�a��Eg^�}��&�˸�n�'���J�����͓<B� $�`U'��AE�7����Ͼ�7�y(Vُ��,E4���ĺ�f
:�S�z��Ɣ���(]��7}��CZ"\��UK�2͚[�\e�C]P�ߖ���}��$���K����RG��j�̹4d�a�.��R�sD�0)���^�
bR��Y56�\<�duä��n�Ao�`o����'��m�Y_�~���rL�F6����UE�'�����2�kS�\�X;N�]3��8t��#��Q=�3H�R�2ۋ� �Dtvk�0�t7��p��R���љ����Ew�W� �qT����"qif���6��*jN�KAܹ�}jf��Bq3��vj^S]v�ì�Y���8���x�1�����I>����8�)9��� X��#���e�O!sQ'������*��EQ�5��r�N# �#%L��R����#w���^�23L��A��*���AZ[W�Q���ٞf�LH��s)P�𵽶�>��.���	��gڇ��5eH�/�L�!
�ͧ�b�耭
��M��0 ��
W�Z:XT���Ӯɐ�:;�򕍒����/ߓx���n�����;�2�*o��W���'�D�w���b���]GEyݬ���	��|�_��!ؠ-��k�yv�z��G�<����	 D<��ې�w��N�}��x���2-nM�Wp����E1�eˑ9r��mb�_�hL�f�$A�tlf�65������9�[�=��E@��H�=d3��f���@����m�$I����OT���|qC�nB+Z�Hq��|=����T� {`Z��+���#�?�ٿ�)z<�[���e�7�n)�,끩�`�2��^E�z�F����B�+�����й���n,�K���g٠c��GV(p��At7�f��r(�'Q���jr���u'1���P�1����y���x�	����t��G9�.���7����\�~�L��r�c�J��b���e�ի��3�eR�|zsn�6Y���g¶y����A��"-��u�P�҄���5��Ó�<k���M��s���^j�D�ܥ)�����*dԱ� O>i	�U��q��㯡�ˈ����U҂i5Y�rX9��t�q����s�t���܈\_+6f�`�$��֤Hk����ӾQ{j!5��Eұe�ۆ�H�#)�Ow{B⒇�ʬ/�����nG��Ӏ��ҭ�*c��C�@i�.t�yf�7��E��fM7-N"���%�2�],�7r}?�SC)�,|i����q�H��IE/��^��l����ׅv-�G��6��/`��<⏖m�>�{�+76]qUt�jd]�&P��X���.�v�a���6��+�"%��`���.�DX+�[�V��-Kl$��`J���f�b �So]�;{Iܠ��)hX�