��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{hi��7	G�����|��4/���YEs��Q��H�9e���ϒ��(��t�.�?�ѩ<�Փ�<�Evj���T�����B�ݰ7� ػ�3��p�����D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[���۰/Zu�(�l�N
nk�����'��m�n�뛗�mF�觴��F���(�wNE)�U��i�ع�MyS���#7���g�/ AXW�,D8lɗ��+�")��p���I��9zg�ڴa���v��QJf������99�}<Z�]4�\*~?���|EL��gn6Z 8��8b�s��d��~�n6�9_ H�u�,B���b��,k�Ծv���0��5�Z?+/~8:�L��`L6����FA�3��PgՄ0�)��F����QuP�����I�<�f��Z�t"�X��T��f���+�>agB�	;� �:z���g�Ĺ�4핤V<���T���5��DxFҘ���zN�E�|�(;j�n�]n�ZV�Zbn��������wxMY�i�C�.dRzC��R��o���H&�,���<�9�W�)6��:YB�a����%~8�ɖ���q �����߮� �[��/�9kڛ�\���V�$���=�}q%`H�*8\s�U7xnH.@�r�%��C=�Q;1�p��&U�����%���|�$�v)p�'d���bmęi�/�PLV��ԟ�!�=�:XV�&_p-�2�˔��$��P��ne�a�dQХ��/�RB�u�m�
9���dM��6(I�0��7��1opm��f�����}�Kv�'����7��hF]5��$jˍ���-�"�Pޏ	�$2^�>_G�U���Y����3=���?b��$�w���Σ�3�;t]���6G�m��/;aP!�_�K;0�|��e���:V��,�ΈG
̥!]/Wn���<��H�jeƽ8+���g�4��Uv�>�����ͫ��Z�W�7�,>/��e0�k��^/������݊�G�����cA��i��.�R����f�3l��T3�\�"ˇ��E��D�P΍�!�L�My�0���!���R����ɲ��F�8Vs�(���^�X�O�i����\o<�e%~,m0����HZ�f�>�
l9����k㺹*�%Ef�l��vk[������<g�2�7�=q߶:�J\^���z>3��<d�� m��P��u���<l5�h
�"+i"1�@T���d��*gZ����i���5��$�#���yx%����X�L�l8D��~.��^����j��$��/7�RɂksײѶo��a�uZΌ_�-�x���@`fH����f�"MSmظ`g����XU�����.���]�Q(��AȌ�Q1�>�PBd�$&x�(n�P�$�w>a���	��3�Kʯ��Ư*�*T����\����I�n��V��,n-���+5��M٫aK�����!8��nxm�`O�9�)��>n���_I]*��3HyR��`�R��Ѫ��f��Ȋ".���ɴOJ�I3Z��U��"|��r�;z�?S���A� �!��.�)G���V�W�Oڲ���EY}Ò��.���|WF@L،����4������޴6Y��t2�G���y�B�x-��aT+�$�����f�p��)���1�!�B�r�?���$M�;�����PqJ1Ì�Dzr��K��&���u����d��f��BxJ�Z5�Óҥ���@��
-Ӏ�/��'���\�� 90ش�����:c�r!�D+�$�N�x��bC>y�����l%�|Z��-�6�)�j�<^�`P�s�&Ἶ��~�2���=��I�{|�̧�?af\C�F�	�(�j�H�F�������e��:w"~�B�wQ���>��׍�	����tqf����E�3��,�:�u�; �3�Yt��d4���=GR�ͦ e���SE�^�w��$e.X�� d��4�
�>�=���O��V�7���vW"Cza��:��q���k��g�$/�V%1@y+�Q��;��������P�'R��9��7��ǭvF��f���yV�����]���A�Ȗ��ԑ�_�����
��焉�
@�|�v���C^��^�y��šZR<|�v7
���g�Z�ȑt;��$���l��:]��_�޾�����^�s��0:!z$�Z�|lhۗ Q�$�Ӌ!`�Kv��@P�)�b�?��NƉ����WV]���4�����K��H��nT���&{'p�&��ý(-k�#���-ν�Q�#-eG�7�x��#�Dt�q�1
�]���5�j}k]�����}<��<��gbb�jZ�*�K�� ��AQO����� w7"w��`Tޖ�����M�Cz	"	CH�
��C��5ݗ<�c������ч�4��>`��.ԯ{���̤N�^�J��Z��0�>`Gi��vq�J��:�[#.��V[��	ѭ@1�oq�|)����]	Q��UC�Υ�[ }�m|�1��}ɻ�Qd�V�����4�G11���_���$H��Za�0̺����� ��â� Y�.=���B1�^�3��	1��귶Q�� rԉ����˼��՜��4ت}��I|���ᩰa�(�׏�{k���� �����#޾1X���/��Cz][E\��K}u��:�q1O	Rko�&bH�����#�֪U]�8٘f����L@�q�l�� ��5�=��s�J��`4[U���Z��AQ�P�`E��gJ��7�ǲ��g�.�^k������'�N��x�[=�B'�op��YL�C[��HG4��1�q�C���� ��?Ĵ8�g�4�.�b�8�`i7n��k�H��PZNL�_yc�#���5����#��i"���Ü(�B�4�L��%������3�� �� wJ��D57P��>��[�ۺ���3H������s��"�!����uW�@T��S�/��x�FOpV�h�4�Y�<����7���pzQ�#�Б���	
}�{�R��v�Ŧ�����Bm��v���ä
�3����:�P�c-���[��Ay`/��Wg����:l*&���P���NEq/���~@�mfb��˽+_SV���2����)oG���!HJ�&:�9���L�`:��ws$���s�Z���Nn�FA|~ec�Gh�@Q�Vg�}K��ڌ
à���WFh��-X�ރ��	kv�����`�S�Xq%em\y�F�
p ��.�a��������n��~�*��\}ݓ~pb˅�K����c�$����F]~�Mw�	�&H{������"��/��0�8�N�1ӿS�hX��׀�.�Ȭm�,��	����%��M�'�Q˘hdo��{��n��4|x�$:��#͆�TS��	����ObC�vCˡ+�\=�&y�Z$����$9�M?h�ڛW8މ��;���>W���>��܇��dݠBB�v�M��|�﬒���O,����	��E�G���2b#h�ޗ��ye��}�d�V8���)[Samh|��Z��,�R�7w�`�%J]���K����7�'�ğ����/�r�<�܄�x[W�g�J�=B�:(�db��D;��No�}�IjU������n:u$Qn��*T�$w�3�(D�����QG�!L����#��6ZhD�I��|l��T�붢ފ�� �����u�������-x���p�x�;���:q���S�Kě`�#*$��ݡM6+�6���Mm�S�V��W����7�H�6f�ܑ��Mq�GORu��T:�~re������L1`���^�Y΂[��/{h����D\W(��֢���w�l�Α�8P4��ᴲǠ�܄���d���:��g�*}��<��Q,��q1<Gu�-|q:�Q�2^;����%%�V"x��;��}����~�0�)"N�j�u�U�8�[U��F,��@Ƭ=�EԧⳊe�����q�/�>�>	5z0�G�Z'H4y�0���-=�0��A�gw�"~����D�ӈ��4tS�2
X{5d.�f��h��QY�����C^)�1W~e����)%����N\�י�>�j>X�leG�ir%�K��Oy� ��g��,?��� IiN��:�����	�,�.3��	l��<�q�h׳e�G��bg�E�8T{�-/�̿��c� �[u����^q���/�����K1ʬs)h��uσ�t%X��e���d�E�3���9���|��Q�o"��K�jKI1���������U�uZE��n��+$�[\��Y���&~2���F:��f81	��QڲoO���[�T�/���t����R���'�*F���わ�X;���Kl�c���:�0w3�C=6�S�]���ڿM���
�Fo(�����x��Q4�E2�({��L��	쮺ӭ}��0��߆,��o�3Y�C8���P
���?�e�m�Z{=r3F4�?��Y�Ŵ!��]K�a�@$aw`�{� L�[CU?�w�K�J�Xȟ�fk@)�Q�s�R������w�ۖ:���f� �Ps� ���ܨ��C�`�dXܢ+9KAZ>��@/-��J��y&�W�j����XDӋ͔)JU�m	�*���[����Lt�VYWhU�o"������\k$inCe8�/��aq�e��٧��)	׻<��N>�U�D�^�K�*B���Y,��ZQ�Z�\��+3�$�.>v�-U(�6��zv���'QTEYc�Ɨ"t����A�Zv�WD}~{���*Ȗ�\����s��������R-}��Y4��<�x;��{�)�Rꬄv�觸$���2$�lRD���3�ZI	I\��3h��E?�*p�1�y�}���yzT�����>)���6l��\%�h���G���S:�W��t�r�E]?!P�/�kf��#3���$0$��"\�M��lC����*�Ի�]ư�oЀ�հ�e��c!bI��ѿBU�67�g1(G�S�����0�A�I�H�Qk7V��*C�c���\���̮7[�<�P��ӫ����jMZ%��${-gd�k`���̪�*�M��>��fc�\D��g�E�J���߹X�P ��L�o�iz��I@h<2�~@e+n=B	�燜@7Kk����H>����7��0�u(vhl��?y�;�K��J7^���%���zo�l��?T~9\ܤ���EZV��β�1z=���G��L����!� 0q꧋��J�O~Ӽ0�/6���V�<4�wgkU�c[vE����"�y�޳�Np��>^"Ebsܫυ���������}���+\^uj�Q�O-���f���hOT�ڀ<�1�A�"�q���rh �J�?�����#pRp9!	��vש�JĦ���������Ǻ� �/н;n�y�;�O�L���/+?����>��F�^N�/�*��*�;�$6�Fp{�;����m*�'���K�	��if��F;���Ն�3�(���	Ay�Ld�������ԇtJ�,y�j��C�I|�+�q`s^����a����w�������WU�#P�Qk!c�?p �ɷ�Zm�" ��l9���-�Y[��SWY��Vk����0���i�[���� ̠B��ˊ6���� 0{�X!9�v�n�ׯ 7a|�$���<�,�~�t|�k��Hz�}��wX͚��8V���{�?�*�g��0^�"\��M���=ɳTr���T�N?��+�l�o/+���7�����zf������Q���$�̜�9�m�%H�� ��L�~B��C��E�<�0�H)G�;��5MXEmtKG"�����t7A[�{��^⏋�x�,�DC�p5�����|�����"��'O��c M1.�)
�OM���o�����F���� �1�w��b7.�ԇ�'9.i�c֫�|��2�E��D�T`��D|�wУ���m�E��ύ �:*� ���E��mw@hlr�9-�\�rC���W��\�� �2�&���`1��SP�Y�+`|)�.ُ9Ӛ`c�U'��7htSY��$�A�Ŕ� ����+��w��)�%@�V�e�F���[��<
L���\��Yُ���FFW�Î�lʵx��.�3�C�M��V)�
.{��$�i���|6����-��J��Z)�ǀ�1xb��
��.?�i���+&�i8�u�a�*������{˟k�y3�xA��"HەZ�$�ТZ+�\���/�8���%jgT��ryQ�y��{V$���)����CANa�|����[A}5���LpW��Q�1�u�T��'*
�)�W���܀�mP�J�������<�:.�CE��![%�����8���B����ϔ��8x{��X��!C��u�+>嘘҈xR7��/�{f�����Ǝ���<�&�K)|ߐO��i�� ���0����T��i�}�m�{Φ��NV�F"�9B�h��i�'[�/�d)�b�6C�O��s����!@�.�xP�÷3�b��/ސ큔������l�A�	��n�K�++��IB���؉�Y����Z���K��tG�����%�m�����g(�@�Wl�@�V��1|��#����"]���.�Oe	\.ȥ�����޶1BI���	��=qn&�3o%U�����̅���-6W0a"&���E� �D|��X�������D2<]�����YA��>��G?i&�wꄗ ]�p������#Ke��K�Ni�vti�2\�7v�.��Y�p�p�o�F���2�>qS���^�"��4��rK�m�
w�,I?���A-jV�$u{�ٸ�۽F,c�����L?��ǉ��e���O_%���r՟is>9G03�����
ᶠ���Q�NA��+X�uv��T`g�\r��h�g���J%^��0�3�1̃k��'����6�?�Gq=��q'�C]���.n�H�_�>���֙e6B2�uxa�u�"�<|P*�:+��V�Q�5�Z�_,�C���p!祙��z��ًnκA����eG�Ie�P�b�U���t�'��j�\#
��ֈ�,$�ͼ���%����^�������yR`�6$��C��i-B�r����ĦJ"�'!�J~��^vT�B*�&iZ���9�����`��H��~O���f3�^�M҃�\[4��ᦛ�WJ�q�{���$�ҮEo�r``ed�X�n0�����8u�n6K
&������m�(W;u1�u���˻�(��0E�u�P_���B��Ɨa
�u�I<ǾB�`�F#D�Sg./��6~�8�AZV�BV���R~/�r��g,�ހ����e�����-yfl��L;��o0��
�� �L����%�6ߵ�L������m� ��y���ݽ����XE�'�J�>���I�Cz��,��96L��P�e7���V~��*�q��	U�I�G���M��V�.�2������H�:���B	��mN(&9��t�����9E�]d=��fCp�IV8�����-a�� ��!54S�y���P��<�n��U�B�_�] ��荟�?N���ăVi ~G�O��eU�������Gp��F;3�AD�/��B�Ma��N�֌e!�d�F`b���Q���P�fE����%M6z$/Q�}$��`,X���h�ch}�j@S�B*��"\g�V��߽�c���O�sn���펁���C^&s�Ů�~��+��f���a�F�o8��$.�=Q��`��U<?M{Y�g���~0h�V[d1 �B���`a*��&�(Y_����o�$�NM��I�e�����a=_���0�	]�!�=1h��yғ�jF'�;��KW�f�mz��@sG�]��Gb��L�N�i6��3@�6_
���k��*.��uL�i~�w7F` ��v����O'��:��L��{R���$������ޓ��d��K��p�!0�>d��I�K�K�`V#p����]�^UBCG@`=������@��I�,�4ږ�Q�rN��_�pX�k�z�l��s�K���S=�_��%HLI+�P�)��;�)ӻ���`kĪ'����-+�ZmXę���qp+޼A�Xy��CE�!MQ` m2����)wt�z$+�� �q�A� Ր)TU�J����*2�u��?���e�{h�IL���� },*z��XՆZ
S�T�"���|��K�/���81ue2��y�D� ��u����U(1"\�S�H��(P�<���p�IH��M�������rj�_&�rw���.T�����d�5s���خ���z4t�㝹� �����אD΢�� :�����d���4�<�o�s�5�M��L�H��K� �dZ�
+�f����g��8zDS����oR�%�5~�U���lD�D,�-����ȱ��L�,�E��B	��Z�m�C�]�O^D�ʕX�T��π_7��s`�
4�l�����[�'��wB�{ɍX���;f�'�]l�4!ڗ�o�9S�h"���K�f�J`�&ʉE���X�O������Kw�W���������çɩHL�c���KB���W�0��vO�����)@��x���d+���^qL���(o��z�"�W�g�{pSB����q�<5�#s���N:V��|����^�P/����/�V�̨��vK�x#'cS|��j��.�{M]��<4�z�A}w� ��Y���b��l�-k�)��Ζ�u����?PCh�uC��G�r�G:�������1�yF�2A������Yl�N��KJ���1w��2�?7�^1���Z|��4�-#�*��*��)�g_Y�gٰFݩ�xs_c"�W�>�O���ףy|�)Q!t��P����1p�i}���ԂE芉��o�0#��˯��A�
��?y���~��T�|<p���&����:%��,.����!G�/I14�����^ՙ4J��]hi�s8P>��P���r�G�����i�A/Zh�,H�����m Nu�t�*�ҥ�Q�j�+�t�NW�Akv�և���v��*�ka��6`2 �Ϡ�*DI1� El��{ǖl@����o�f�<&�X���n5V$�?}o��>��S܋Ϧ�����G����2���K�zf�n���\����oC��6�Wڢ=k0S+D3'�0�+���e��C�0�9>��oǅ\/aC&eж	K b���D)����2ٱ��R%���C���0��sT�[�n�{wn7:G���9j��S�:\�9�ؑ}�>'JYܯ��ܞI5��L��aa~��\����M��3�Q�A)RB�j��;N�e�m���T��n°Xo�4��7�u����5�Z�q�&NI�up��c}��=(ʨ���G#��"�%�c�C��^F\б6��7:�ǣ�@*��
�y=���	�@Br�#��Vʛ�?�i�*b2&���
�,úy�3�z���M�."�>O��b�<�:�M�.N�'F��.$�]�R��^m�Z��[(�
���8,ܧ��}�ɟ�T���%�I�[��q�1���آ�%u��1�����S��e�݌���K�[�$�m���Ou�XF�2<�{�S�ͻE�i�Xm�6|�R!�p�34��p��E��1�&푠$���k�7�1�*{�-��~*�*�S��-D����+t��^�#`�i�ղA�(ӟ��6��&LIr�o��<�T�ӓͥ|lf��ɤ,�����!rZ�`\)�$�{�K�.�ς*��s�Փ�kq��&���V� ��t��=z#��_m��m���,�^�"��c���_�DaUN��[s~*�8���:�↑�ʑgX��4�I����g*ܹ�V�O��IP��/�:,[;��zx詮��	O��I�˅��iO�Z�$�Ve�v��J{�ϸ[Ɲ�2��W�ң�}�ݠ$y�1��������s����P�.������9���O�
$�ʕ�b��s616~YC���|1�:�����j�O ۈ�{oQ캖��5��<���n}s���TU�W$��y�if�b+�J]ɇ�1�J8"d�]�W���OFM�H�.P\��9�/ǭg`�pYD����^\WY��|��L�V���O�x�����$�p�K:��8=&5I5��Z��4�E"��r�
vP��J��g��k=�Z������ ���3�Gd����P��7��#�͝�$��u��81���d"�d{Ç.���Q\��ڪ+�xA��w�iFO�Seh�`#��,[lm^���X����7i;N_��)Z�2��Is̐LS��g�Z;��/�S� Bo�2-'l�#gl;��`+w��b�{%Z���*�B��%���
�6�F�F��̡�cOL+�ܑD(.��$d2ɶ����� ̈́ŀ��R�X���Ӆ��BkU���T�.[��"�朆��o �T�m
Ņ���U�I�k����N�6�1z�Ff<r�B�nXCڡ[�J�q��B}(���s�t'!�{Vȑ�] 34Jb�&uU�o��5��b��r�t�,.4��t�ڃD���i�2�V�Y�E
Jg;3�x#x�
�=Dq�W��={Q76y/�N���O�(�����*�F�w���!8@KqGe������'˼�]z�4����c^M�@��E��&�c��mԑ�������+����s��cG���K�|3�u6W���_�)�<��빲%aE��D*�v@��l��-�t����^��0�eγt���=��VAT�F��4��h�PPYKA�_u;3�D��tƚ?5M�NC��5�������GP��ߛ9��g#��z�تO"��&n��J� ����A>֨Q�2v�CZ�s��/z�MN�[BE�vC�3�m��Y��Q0W����h���ced���q[�����5�ԣIƸ�H����CgV�o�&�����uh>����`͵�'����i·��2�ʡ%��๾��R�"�γR�Ak�mt���.�_��SxN�Ȣ�p%&*;�hnu�R~�8^�P��U�'�xs��1����C*�2u��_nB8�6��T�2�B��Ѣ���1�������P>�,��;zE2IS,'��\��X�編ζ��}����G��"�*X�V�:|�t�		�E���X�<Ǹ��Ö��:�����w؁���H�o�f֧�xuT��i��(�jtE��	\�5�qR�]>�|��B�o�ҋ�W�׏���KZ)	>��q�~��o�mK�m�ݙ�Вk;�g��p�K�l�(��[>��ȩ!�c^�pF���&L� ��|Sԣ ���OW��4;�1�����̥(�{s/^fi��{(�+�'�r��=��d�QK�B��������\ۣ3v�^@��1��+������P��r�G�zR�<"�N-��)A�7�pÛ����"pAD���|v�Q8��oHi�`�����d�vCjG����G{Ck��d6gV*��wg���m������60Ab bgV�2���7S+n����� n{8<�:�)Qﮕ��$|�C,+8Q���M���^7�F.l��>�'f����o0y�lH�; Q��<z��6ɸ�/�w-u�J{�ZL�N[W�FG���y&� g�xr:;q�o���:��5�	Q�1#q��9�����؋T��=��<�Bh�I���{�~�9�#α������k�Jf%.�め��d�;�5�e�����5���4�C�^��0�� �*ܴ.%y�Qjq �J��������[��jA��V�.�`��_9F�g�q�v`E�ƾ��O@	�SX�l�`x�'h� ��FÇ�/&�׾46�s܈�}�]��7�u�NUsG���P�9��n�n���^�ۼ���/�uM�������֟㟪4Mǽ$p*ͥ�C��Kʸ�m�I�f\��VV+�G�v7�-hT����3ݠ T$�q")���ҷ��r�3�Y� ���Z#f��9u��i;�^�+�R.k6�$:	ezDD����4Z$?�Sq׽^�x�Z���A�j�yL��D2-�ot���&�{[�B��;y_N'j7��
�u'��l�q=�Q�����8�����j�/4rϙ	}wת��)^霏VQ+D؁�n�T���K��ҽ�G-��_����M�d�Fv���sG�1�J�1?�wm���<X��N5v�7�C�Cc�ğ��Ya �%R���J�E.�A��짥M3�/�Edu����s����M�K��%���Ga�%g�8#��6���8V�f��¯�?��U3#('�E+c�GVP��b�Xד�U��t/��e {���-�V�#N� �O�y�ƱW1��@��6��\����,'�m=���Nݐ��xw���PW����c�ӝ����ac[�-��n+摼n�_Z�+xݥ����n��p��ދ����M�;(Flή{E��]�vkY�u�爕@��)~�-{�q��2Pܘ����
e~1�$槿�YVr9K��JƂ��.y��a|�~�R�'-���X ��|�i��t�����$MdQ�z��<&�G���|ݚo��u)=ʩ����d��-\�+tG`�ZJ����.���.�)���sRպs��-Ƅ��a-#-�;�P������(z�� ���\�&�1Q?r��r�5��c>���]�����㘪�F����|W�b� ��f�`;���ޠ�4�d�FJ���l� Ru2�W5{��<K�Ŷ�8P6.����0c����wcp�v��#�߅j�lglq�Mt@P7�:��0<m.C�צ(�^�s��r��F>�PcRa����L 劖|�i�N��y׬��M?֌F��uR������ɺ%r��P�0�+��bw�/hd#�+e}�1��в��Z�I�/���M=�F�	�o�jcl���Z����+jݧk�m�9Y"�-�4Gg�2��W����pj�x{��x�t;�x���k!z�M�e;]N�I�/�H΢N<~�u��s]�$iTF9�;ow���5ޥi]P\���yG��AP%�%S�rb�S�i�K���W���y��}	��
}�'Xhs=��:�����UR��7�&@<q�/����>仍�M0���=��"��P�O2�'q��k[E/e�B��)��-c�t����7�-_Ch��LC�u��M�5�L��>Ma�\���
p]˅�=���� |��f	eV�I=�Q�e(���� �3����
�O�w����I����E��r�AK�̼m��!c�'���g�b�~y��j��}�XP�tnD��0˰��0=�S�u5Jx�K��F�T���J!��wu}��چ;�����X<��wf'��>n7{XB�Ը4���^!Zh�:�Y{"4�'�j�Mao�GB�eE��/�jg'�5����U����Z�	.�o��Kz#�74{�������x�����)K�z���	`���`���I��3�PO-n�������ՖzN���hrk,<�sP.�Z5��+/��cҽ��ƶS�s.��e�vd��\ #�v�^S��嗂��a��p�O�n�\-��7�P0�1���
����R���X�7�7fp���c�+|C��3��t̉{�mW+��՟D3]I�>�`�g�m���xu��ȣ|o�,�(���K�l���ӯ�g}�j��qlI�E�r���b'���Z(��%&*��C��������A��c>.���DI�������8i��q�U�*�|K��OO^yW���Up��s�r��k��O|�:�_��`@~��8��9� �+%�qי�G���;5�h�w�-���F�i�f�b��v!�z��v��H%�u���&�]��Қ�W��w���AE,�BW���QE>/I��R�?�/׬���F��Rc�֒<�)ξ��I��RV�>Iտ��{%���5t��a��rh}�A]�d��!�Je7B/KU�O���ze!�[1O͕ӧ�^CE�~&x`�hg���}	^!���6���,tl���R_�qbo�Py����	t���qIZv��"�H���
�G`��U�tċ��������m��%�b�t���*�������[�:e���ë�R|U�ךZ�k!�B&y�~����櫌��
��R��.Gҥ���;v����Z�}�T���Z&wV�D�)j��v�f�kj�0�y�Ř�dtbՋ��+�����Iˑ�/PTv�2\����S��R����� �T_���k��SXEp3ۚ<��֑P��#/�cO����i����cqv���!�t�Uݭ?�a�� �(�#_���l��]mi|�1�%�Je$�+�)�pQ�Bw\	��|���l���9�����DoT � n�6ʞ
�0�Sf���18��a�i؅oZ�b/�b��E,j��L�[/���
�c�q����<zH���e�In��Z��ݔd
�Hu�ٙ:�l}ty��<�U��LQg�|, �ڬ�h�S��'S|FP�6I�������՞2.�uu$��\��o�a�5���޿2]1W\����@���A9@�y�@:������}w�%t��bDcC	�k��H��δEx�rQH1Y��������]>*(�;즨��2tz��o.�#��fȼ�� ��HF �����׻��(?�B�<�>�m���xQ��]#o��;��߈'n�t��'BD���Cm�
�����[��8a.r�|���2k�䭝����
Z:�'�6'K��u
Jn�[��j��6�>da	
zX'�R�c�tŁk�brd���%��e����C��.6��P-@��l�A��x��B]����ԣ6�F���s�7�Jb:��{Gʀ$�o�u�x��D�%I?�0ÎJZ&`� %�Ɍ3:��<[����L��p���2�l��9@�۷� ������{��)],W�ǛJ����P,ȸ�x�{��J��Coc���5}��$�B�W�[��׃��BJVFY��9\���.v�.���k�e{&�1f��!�o��A^+ײ�+�[�l�9�.�w�&Z�����ڇo��l?�Wuݰ���������\��e���jӇ}�ER�,h3yFS-�iu\0��o�|�'��_���*X�V���{���s|K^����y�2P�C���2�mT����z��M��\(x��n*��:���G��!��]���ω�,v��"��.������8���9)��|: CU�T�!�R�=uE��2���%�;=DU��ZW4k�Du�~�	m�B�wu_��[
ժ�����q��I|_a:��-B^��ވ��rƊ�t��d�?��%�g��Y8���t��Jdd�s�ɫi��hc�(n��]�&?����ɓg5�T	� �r+�.��AJw���)ً�z�Ŭ"N����x����(8���Bحٌ������}�̳�#�6a��X��ۍm}[��l�8���p'5�U�F�؀�Tߍ�;��R�?�G��=n�#O�d+|�II&��Q����ȅ{�����ȗ.�X�����[8_���a䊛��A�9����+���&�tC��u2]'�lX���W�O��o�u�p�Z�	���x�[��?��h���é��9�����<c|R�؟'12ۃ����ɱ�;�ɕ8��~h�����i���2�d�	-f����[g���;��3^Z�o�A�ꔈ�/�(�]I���P&�:�"Xf[:���\�����p��B}��X������� �q���]��/��N�|FL��������e�'r���+͎�动��B���!}�c=o?l��I���D�[�1�}0,E�
EU�i�o207��֢$�˙B�m(_���glQ_�P#aFe���գ�Z�\:�@W��k�$������
Ki���׺�UW�|����:�~/�lɿߝ�g� //��$������_^�T�� Ͼ%�w�i{a���$�{z�r�c���E߂�W*jL4̔��g�2�x,5R`��X��(�q����O{\?&OޜorN�w;,^�KGJ��2�L8�.y�/���b�\���%;��?� �R!u(���e^\��є�<V�v>_3�5�`��mC��u��9k�<����+���|ԣk]V�c��}RR"��,Ȧ�����D&n��H���4D!-�	���9Z�r�N&�$Wr<&j��nGӣQ�jW�+1mq�J��(��Qɦ9�O���Ra��9��}L�-(L�;H�c���6"�O��H>0���l��Z��J�L���t�v��z�V�y�t���Ta��*�d����yv��E3�%������y���=3u"���MK�'���ۛ�:;&���H;rc�|�ϛ9p�+Ν��_�Ho��Y�a�8`��������WאX��P�}�� ��8"d�JS:����Pj�Ƚ��iQ��=���R�py��R��F���K)[���@�H-PO��8o�`���D�0Od&@��7>�H����$�qW����V������Gf�myL5��2�4�1�sc 6YJ��������@pS���3Z?M���>$�P��5��Sg;1���˖����=����ktN_��=aß�ק�n��	K�K�%��.yh���"��]�w:�5S�36���98��"Z����G*c��U��;a�&/�8���+�	/�ő�̐*/`��8;���=�x��r���\`)���?�5�*I�;*ג��%���N��B�/K��o���N��H$�ۚ�������|������x���=��;��?	Z0�jj��Yо)i"`I�����Y ���Ǉ����`��k6���ԉ#�*��̗W�`~^�hF�~w�
��$km�ky�K���c���`r"�$8�!�I/��,�9wE�q�o[�錉�M���a�$nH�y9�r꣏8P+v@؃�i�р��W�,���:
�k(P~_��L	����Vh>�����P�����z����6�@�V8)�����2�F}���x�>�L��"Bg�:������A	]���MȮK-�ƳE+ 
D�{H짞K�8T�7�൳�_�*��(����I4kxW�uan�/q�Q�(��w�%�����ê9�̓�֍^V7��N��A�b�a������B�#j�ӽ�� ��dt�KUb��쳻�E_����;v"ߞ�X�IY��u�~>��`(�l�?�:�ܓ%�!�*���Y���2����W��\�R�$񵉤� �^��2�i�ȷ)���v��:�Q�tjw{�=�����l8���	��������͎���H{`�]���]�g�?b�-\���6Gs�Z�:-����<����W`���p�b/qN�'-�Y�X������I���k�,Ќ�=�c�dh*v?��z�֣�Up'�t��S�FS `�E���HJO��־�&�c���J|�Y��<�"R#Y _�~QN�Z�!��Q@$�i�Qf��@�gn�j�}�͝�
@x`�F\����P��Ɖ���;m3(P^�b���7`�omÔ	�WB�7�t��U{>�Bd�< j�qh1�ݒ[:CE���}!��%������tǉ���%�S�g	m:@�Z��%&mCf=͙�MU����1�w��y�=�6��Ss��P�Ʋ��9-�����g�&�x���wɣS;tu_���V�r���qig�^{�c9���G�ҷ��dM].�+u�P��Ct���'W�����l_@��^������nO�^�ȱ����up�m�������A�<�_�u��F�zV����@������0�����+j���¿&x���hb
�#�^��9zy����>h.��l��-�:��mJ9�3ғ+%��,	zR�q�\�r1�Pt���bd�˫
��r
 vv��lH��;ü��wb=������	r'~`a��-������-#�v\�w�ޗ���V.o@�J���f{5#��[H���s�zP��0/�#sޓ����r9�:�tҟ>�5��J��}�6����5�ZVVzAx��Į����ϭ�$s�� ;0�q ���C)�31^V��*�	`rX�K���KT�S.GuP|$�� �r���+�v�m.z�;w�Sa�B: (���V�l���7�7��$�]Hp]�Drsl�U��E�����E]1���z��+Hw�z{J5s�ݖL�5�։3���u�T�������'�"���^���ʚ��u#����F�l{g��y?��K&���
7G6=����Xv�X���kQ��Jx��uT�0����~�����
�Af�S�hBO��99�Z�Uli�=�r����չ�?�yk*N�˅�w�]�	���C	7+tM�S(�P��O�l����W>��LA#Np�xB��Ph�Y�<6���'bNS���KD�x��%X��'4���0睏5%X�&"ѨX�ST�N~�o�Ry�����?$�D"��d���]�=4��j� UP�]_�I�!��QJ��9�3e���\]*�c�N���)�mv-8~�I�v��2����S���&S���q��/y�kv[s���TE��iFї8{�Q�y��k1�~�k�ķ��԰y�.��	M��9�O����3��Ai+��"1�B�q%��\x�m�Ԝ���F/�ӯS�O#ʵ$2{­D?��ŧ[��!f��*]��R7W��B�S�����-)�,<o�'�qd��1#��[s�a���ؠ�X��9Ks@r���6Q�����&o9Z�2�p��O�ʻ�#��,I����%ܺ��O@�)PBz� b\<��� 3���\[����1O�n�%��ja�k�	ʶ���z��\
Wd����m�������=q��T[��qD�1;k8,1!��bOή�W Q���<Z,�L?�(�&~�QJ�ߵf������ ���s�Y��}J�^��4wWk�_���j�UEW���PD&��uR�v��A�v��!\�Qz���ؿ�^�ZK|�ęU�;�P[�#UB��3b���kka %n!ά�cM�|�"_�"�(͊p�_���}�R�6�o[�.V��)a~���8b@�ƟPи�d���VO̴t�M0ݣ �n�Fxn���@��tɧ��I*,$���l�
I� �Ү8#𫴬���\��:I*�_I }ݪҥ�kk����Ƶ�������c/.� kD�� w�ۤ5FC�Կ��z��U�'�y],8_.+iS�.ȩml�e���j�������
K�?�>~���;����ǘg��1x� (2�.��[㕯�{(�Q,��F7b:�4WϺ
�X5£�E�z�'uW]}���H,�P0i��)8�5�5mZ�s�4.h1�oa��Y��j(͔ѩ�t�dEcRwq����S�gKsL�ϙ�Ns�����$����;�&֪;P�J/���H�M�&�)-b�GNA4H^�o�l2�Á���Ԛe��"��J�����˯=�2�8t���zt�h{U�����hm�j�|M��A��:��m��9�`7��X�=��M��[���
,�S�B%�.H�Aܛ��NK�R��N7��<v�Y�L�jSo���흻���u����kφX��'�;��|��\b�H�aU�|�����d����]��FPNZ���3�
�)�V������+���T���,�S#[������pxc<�u��78>���^0������M��JN�2���� �tZi�����Zг^������Q�l��?پHϡ��8�n(�~8�C̨�?\f�1���
l�������$\I�aqz�sYM�����L��D�!_X!%M8*�$D�q�5s@�})�-i��C7r� @TN˂���hP���XY��$18�_\^��o���i��ҚS{BɃ4��J&���*ƸY�Ґ�sUZ_f�r\�����5���X��j&�|��h9�}��9s�N��W�y6��/�	�2*�#�7�)l+��������Mj�I�$�;�ӎ�
V�<�����0����ۯ_p��7�t��`d�D�2�""Biv�q����F�k݆v����%<�\B�j=�?�[`%�y&����{pQ�Z%O�kr4���lȪQ>��4�bnp�*��(X0��/&�r�_��4�=[|�h���Ah�}r�D��X�~�[��!s^���������>���^�eD������aʮ-f5�_�	G%���2�%�P��7��;+� ��ݭ�'X?�4���_PX�w#���a�.[#1��Gh���71�Iqp7O�ݩ;��S����w'ӯ�������656Q\T����V���s�*�T�*��}�i<,���!횇�8۞�!˙k�a���������x=�` }�6v��N7jl�/�D�d�<}`���+dU|3�
\�G�#���я�x��@x��}i,Os�e�FBH�Y2���]-�OG+Z��Ъa���[6贂S��Эd	]�f��<Jω��$X��Ȭ�ŧ��R����8��ǽZ��M�Ƨ4=�S������{H�9�o?T�8j� �
&���_iCw
�F�_!O��<eċħ.KY���s�=7����}�����#��u]��P�:�\lm�{?]�p�8U1�>���z��n�7��_�$�:��������#}��sg� ��C]�l�Q�� ib�gI}'l��j*i�M��n��-���+>ڵ�ة��2�0�t��{��U���Y)#D%�ƒ@ԴA����8���H���#���O�]��:��1>�����^.6{T<�1;h��P�_�y!\�2�[�Ѩ�G�$oI��(MCw.�#���oH-G#ŽY�ʓ�����A,
�r@��˗ؑ�l�V8^�A�t����_�;�@j�%�x�A���+mȥ��ʪg��>�\�˙"cC���X�I���N��:b�ZϮF�
�r0z]t�4(5u'��aD�/3Fp*�n�m��z$E��������Ȅr��G?�E1䖃�4�q���<�RG����`kj�YP|�,\^����^�����3*�tu�4��8�&
�E+DUpY�C�[����#{|��Ţ_[�dט܍8�W�*x<��̺{Y��1����P�|�^�<o_�3���؈���|Ev��g�wQT����廛�ܩm޶�����J�����%�T[��Z � �~���u�R4��
{�4Z.f�ZNJW����?���R�.�y��`�WHJ
�r�i�"�;��u~��*اfd{�)��O��ߚ��b�< Aދ0���1�����-;o�������LM�B�����h���4fTtY]�(�(�ކf����O%7ȥNS,T����)$������G1[�H�����
옞/�	t /����
~* ˩�׋�U��I� ����EG����p���ߖ�q^S��,��&�WQ
�¼�:Q�ו������,R;N��1\ Z��Ͽ�=����wH�N\b���wI����,]��;�E��[|��t����k������nx���F�<�q���RW�B_3�T@�U��3�G���MC��8�Ş&���ٗ�ej����-��m[�^汴�eS]:n=@0��_k;G�t��I��J{-�LW�aT�岐��ةO#�{fVoI�*�a�y흨|��[9�Lל���MW�y��ȗh��Zf�L����2��~(s����So�K "�;e:JaօԂڇ����������]��RҖ�\�^bYm��4@�j�j?x����N'��V�S����1&�9'1BI����!���yC8����S�u�,6����qF����X��ԃ��Z���qPUI���ԫ Vf��ˠ��z����|�v7Ԕ.���}�A��e*o1K:�x�P��v�׫P��כplbj[bNyh��d�hckM���(H����!#��4�]"� ��ƍ�JOsk+��_&���?j�>�L�<��d ��,H\�7�,�/:�����BԄܶ]��6!��a.�=#"��r_���RR��*s銉��%plf�eH3��So����2.J���]z��ϝ#�P��J��i��f_��sx�R;D�� ~�7 �ċgoM/I�,�^42�A�q��	�<�s�|@@:䮑��mť�P�o[�p���2��h9�ƴ�`�$L�ogOb�0g�d<]�Z��1�`�г:Q�m�#?�H���eMFe9>����w��%�*O?��2�r(�9�՚4�;	A"�3`��1��r�?�������ԍ��/����;A��'}ܵ0�"����'��jM��X�Q
X���R�9��$���}��ߩ&���f ���6����DB �a��^�ƺ٢V�`����yk�3�θz���֭j¡����X8r�������&�����Wj`��'�9��W����ͣ?��HMs߆D�F=�X{ݺ��R����ͽT�"~���m)�3#�5��
v��o�h�m�4g�,18��@ON���$�s�_|,S����#U`~�rQ+�������K�Y?$����6�>�Ч�6T��Ǵ�*�"nҐ� #LkeJiwqG!�k�a{2��肛�."��L:�U\���\�7l��I
�,6��f�Rn���U�t�Kz�&ۮ{ݯ��I�o����)s�^7&F�tA=	�Iݓ7����`ѫԎ8E<�g+��X�Fk�ݜ���V��*�8�o��_ו�� �U�AO���!�}�0�i	�/���D��~��.�� ��v�e>��R�*;#�vp�S��0Z�Ώ��Icb7ߚ��P������!���v˕?i��W;��c5�C�Ow��ݪ��Z����M��a[�q����]���A�"?�v@���'
|��X���ޣ��ku��]�]MW�+N���=� �����櫴#��S$��:�����&6��-T���"��+`0���[�S��� ���e8�������4�f�&T;���N*)�as�"���a������ѥw�TJ�:���i�M��)_��C�(�vӅ9�k:CK&�|vx���,7�n�?���ק��M�8�A���BL`y���o����O���e���~��}�����jH@8x�[V.��5�>�L1stASH��x?�c�^�T��W�u: .ju�TP���N`Ys�4͌ �[���S����fr:�4���ϣl��6_v3�	JWyn���ЮAœgT�})?9���������B�Ǧ\�j@�����'�T@r/��AD_◱�c$>��[���L�׵{-|��y��я��*�q���Y����-5���u:yr����gqǂ� l���*}X8�XI_[�O%���@,���s���[�1�Y�=6�R��`�n��`��۠�;���[��:^���%<zu�u��X�pݻ�p�+-�C�����ߑ�	�5��-#]є�w����~uwp��E��ϓ- "��E�h`;{L���p��"��ϗ������{��W��(r�S���mX�ʈ^�8�-��&'�Y>W���榪��I.�(a��&��h��^��5�6�<�ߑ�|DڃRP���J����~�G��E9V���?�D	�еa!V��>��5s�Z��N�"=p�����e�e��,�{@���]1 ��(l�����J�
~��iϝ�=�"_l]W�x�a����!��w�Se�V�:��s�,�%����z���d-O5�M��l?�d'N����̵EaJm�?ֱH�=�dh*���J:�~�(���M�vl��7,z�Φ��}+�(�ɀ���������aS�#��M������v^ǜz�a>#�eF,o�6���`hJ=Q�P�p��IB)�bO�+�G�v4�:G���}���%��N��kNW�eY�e���9�9m-w_�����S~.�ՇǊvH����������!uBm�*¶��5��J�G�|�5�����f$qC�kmП[n��������<� ���#N��=D�w�;��(0���#�E�O,0D���>>�փ悚�+�WC�5�Ս�&�phF��?�JH��TQ���Jd��tq��y:�8&ѡoc5a���c�xÑ����c�x�hARm��sF�zs>��e%E�@�+^ֿ/^�m;�a�E4�T�0�<�K����qBL�n��oXS>�^����C�"L%��ӱ���Ι���ț��/PO{�%z"F6ڱ2�F�W�1N�ٹ�0����@��Fz�Jz��xS"J؊a���J^X��L_�P�K��K�kN��In-,���ϩ��m9��_����Φ�e�^7��$�+�i�"�#�tu����Jk�Z����Y�#N�m����s���I�iH�W�,�$�h��<���.ʢ�f�^�b"�V�.-q�p�#���|%)�Z!�)���/K�ަ�VX��#�]Y�����d��۽����T��I�deIϩ�B��u6To��'��Y��(���b�&����>�;�o�P'-�ž(��W!67�A+�cI���=��m���0��FD1T_7A��0�P�u��4$��J�.�"��7�����ܶϣ"%]q�n�1Gԧv���ں�6-��?л��?)��чPU���SA:�,O=�2�"�lu��V�|�ڼٶ�6!%S|l�Е�iM>��gH�Ǳl'�!zЬʂR��`��8K�V`/�#nCU�$���}�A�zv~�V�PPLO�����D�Ot�{:��4����(p0�ګ�.�W�͏�2�/G�k�gR=�(��'|���)�U�r 7�ly<����ςy�蹪R�y�}^����}���*����C�CLx�8(��*����2�yeB��AU;���s�����߸;t@�2��5�L��>"���d47)�3�0�o�P��*�]XO؝4�t�+ˮ�>������wA��
#��y�vs}j(��V��$�ezf�\����P ZM6�bZ�.��Ռ*S��vv��O�ȉ�q� ����s��fd'��8:d���M ���كxw���S�C:ҏHW*���ִ���լ��ڍ�(�.�޴�Ա-����7Qr��i�؀2p�3t����@J��J	���j��<9u�?�m�\�K	<h@-S)P��w��(��̉�Q���ؼ&O�5)Z/`��ԩ�S�[����3���&Z�tŐ�o]�a+�T���c��q��@�������@���ن�Rce;G�O�!Q	�I�j�I��E�\?��(�H��o����a$�R0�2�q��%���,���0��ܓ�H`(�9���n=y�,�MCN�+�G~�u��mq`��@��;@�
5�C�F�W�`+q�؞�d�-���5�%O�'��rj�e��d~����I�O�ͯA�<�
�f���q� �y��QN���G@�����u�8@��
�Y+τ �����6_w�n��x
��Fk���NJ#������ ��v�&�VB���0��aD�{�(��CX�a��-��2��+Q7M��y�U�Mg�܂��{W���[[����J���yd��r�/��GAn�/9�P��PW1\U/�e�in��}
��93�n.������]P�)��%ZT�t�{EY|L�d�����z,��3l��z��>i(j}�r�cQ襒�o*��L���ɋ�~��ᔴ��Y}*,;�N�1\���Pxj㣻��Ԏ��oǓ�8�:�k ��U!��6�e
�!^|L��8�֜�Qt�����X��Y���!����@h�"����%�0}M7��ۊgD��]�0�|��U�LH�9�-2P"i��uǨ��hI�R(-�8]~5	X'͝h��ưH����I+��a�se���Hq��ʧ=��!,����æ���ё����{ͭ#�PnHw��߷M
$�	�Ӥ6��Kď�bFI߲��s�l�2�����,�@�8�����.;����!3�y�� }D����Ťq�/�����B��Բ�N�dT��T'�tpq�'uN��W9�d5E;�y_v2IVp�%��W)�Mk;��N�p��i�f`�Q�b��SlGV����V7�
�OU��g�w����Ú@f�F2�9깪�iI�vj�����ڸw�\!�Hۻ�SO�˟�������)�8�oߨ,���-���^�z��z���p����M/,X_ ��!���U.TjC�)7�q�
2��gy$)X*b~����(�q[���|q _�+U��Ѧ}w{Q�g4x#ϣ6WI�<�w	
x���Nf�}r��-n(��x�v�mI�$p}��E&"eV0&�A?�"mϱq�ԶxL������{o�绠��.^���;aV���_��g����Fx�et����s�a�;��e���ֻ楆����u�WQV��h����S�D|�i���~��G�-��H֊��H�\߯l�*�Q����5���Y�_�ޥj�n,B��D4'�����[P+���}Ts:�Ix�b���mX��n�l�T�4��M�����M�gc�:΀���u���-�K'I�)|*�i��QK!^G�M:�|�y���,%#��/X�]�wf1�Ӱ�W���B��ԗ����^F)��)Ɇ�z��O�����Si�r��'�2݆u��	��};6�$�$b� ���q�T�Z��s��Q�a5��㐝���\tM`0p�O�A&�9��z�L�Ϳ��0�
WwzYm�p}�6���
�m�M}#����]��^0�'�7��s8���:aH��6K��-J�^)��>p�j(�|+ )>��jL���{7��o{�o��n'pк�zs�x�O����Հ��p�lX��g��R�l�!?Ѝ ��5}iއi��ۅ�dªu�b_�*����Q�L8��f��Z?'��oe	Ġ�<�X��������Պu)���qwC������[��������ۯ�Ɨ~�F�u�q@����
�zC�yt�K����\�����2�t;v���q�-S~J�9RM	��)	���2��Y�1���ͧ���隼�I�<�o� aZ��н�JԲ﹓VLJHb�Tg�ӁU!_e�b�߽8���#����L�-����5�P�Ȧe1���Vi|-)z�L,�L7��=Qǲ�G�`��J�8}�$]����,Kz��Ŀ�ZN>�L[�/�8�Oa�ߜ�"���5� ��L� ;d�+���BJN���{x�U�-c1�E�7-�(�Bǵ
��5���E�x2	��V�R7Zپ�HܵG��s�X�W�.��cb���z��L�-ź-�9E��E[*?J���sb�*��=�s/��΃,� �lxx��b�w̎J�*�BQћ��k��PK�d�IuV�p�ÛJ5]y���+c��SS�;$�Y��n|��,���P�WD�l��PeG1��G�}63i���ѝ9-vEp,g=]����3n��PI~>O� ���C/�S��Fc	7n`�SҀ��8h�@ԑ{&0��m��>�&��Ф�'MX�nKѩ�=#���)K3U�R�X�fq��0�[��R�X�A��R%��A��a���ou�(��F�9c_Oo��ӧ�9:��g���;Y$_}�3}-�����Їk}��"�)sض�N+0;/�G�eMUh����L�����"f"�5�hc�@��a�^�:����{��p�%��m�Z��H�8��C��\	3�j��ȵZ�s�c[ڂ����@��p�V1f�s9�=~����y����?�L��:��,���;�KO���L�G�x8��S��&�֞���H�PJ�=�دPN�y˷G�A�fB{y��K���x�X���;�#J�MQS_�C��#R�T����w�\���Ӵ���o,���HF�#���I_~���Fj�PW�ԑ�y.)��C`㹎r��VȝJ��������Q��łE�:���m��\$�96>N�ۆ��(u����Y�Y��9� �A��T��/�>�j4X���v{�	��լ06{Ei�`�Ncй�?r�?��w���ƍJ��`n:ʂ�bQ_Z����ëG��+SQx�>|[%Ot���6,�i�pNᓘ��S��%ll87<'�+d1��z	L}c9��U\��-nv �]%�-=}��nh�3[A����F�HU*��(�	�>Ȝ���D�e�+#�ah�0R����B����M�s磼FP�[������y���ם�:��^�f�Uo�qJ6��9�S���A�`�_��0_�^(A���"~!��]h!����.��u ��-P��ޫ�l7�sn�Z_������d��!����#���Wvp�;�ȧ!�����k���_��1:u&����Z�$g�@Rۉ$.�|V4���5�"B$���!MḃJ�PD�5q<H��]������YD��z.̺ʰTI��Fu,MLi�\�E���GV�뤹&��C��-������ՎP�l �����[�ީ��YZ΅
�TI��V�)B���>�V|t'(��\@���¥ ��ܡ��dgŒ���y�&��٢�Hx���/����=-Q��WT��̽��ˑ�z�YB����#et3�W��0�{�O8y����A�"QR����O�:�%��|_��9��ʻ��<�<Gi�<�8�>8� �,��@Z�8d(����@TQ[ʴ�[�cx]�k�εP���p3;�-�Y�9FD�� ���{\f%�6d��N��j��'9�u�SZ}��E�t�s�$�nԢ��UL������9�뼴��`0�Zx��Ƥ���}�|��'Hڝ��6���;�`IoZ�w�~U�.��Y/�"cۚ��}���VP�����"O�O�f�^��aOl��C0�"@֕�w6�L�2F�10Cz��Fܶ_��Je�	�Rf���BM����e�?��pD�5HCz+�q&F����hK�o��z��Uښ��*��H?3�\����/��(�q �P\������Q�z��K0i��W� Ǳq
c�:���c���G��4��2��� �H@�R�T�D� R� 2��:]�y�*]�#��n����muhu�U��WP+��*�:��>�y?CSUJ\����2r��|
S�t&#�
K{Pd�\˟����d��_\�,�uc�ٮ�a�&��kX���ݝ0����>Q���_*n=����$���B������B��e�3
t���!�V���7Dm͘��M��1��[̩q�8�2��ԧ@����5���ɂ�� CVQ���zȧ�qR�5ѸЊltU�,�Vޮ1%� 0��5���3kGC�y�*juTC/��"3��&�@�͑�3
(�P��d ��Y��d�놐����<�/�-�������n^��"�Cʅ\��`J�<G��ɴ<����h�w-�V9�����N�]�X�Kf�)�[�}j��9��˷��x�"��ڀ�1��$���`�(������Z��0#��XV�Ɲ���G�oT����J�~N����'���]�I�yLQT �x�O�~+��Xj�"�]���k�͢�9�0�J&��{�����q��E`���~�A yY���ke��$�Ъx��J�V�Vk5�kv�2��<�O�t�X�&�iZ�� "ǋ�v"b�����sQ�]:�a���	"��nX�2��2�6C�MW���>N63�IS4"����e5�[Y��J���r��F�W��Il#����,0as?[V�M�ݻ��N��͍�Uc����Qܨ�W���wX���St�{�ީ���ۀ $��!@���/pn�;%�I�%��\��	~E���0�Lڲ��y#���gHo�?��TY�@&���е�'9�{NL����� ]N˸z�����q�#�#Sw���IS��g1���;�9SI�`�#a:v�:X;m�y�sI�r�4�itLV�~��b����
�>�ąGm;���u\�.����*k� z�CT�G��NiRZ�F>�#�B�N�J&����7+2�3���R��5���i�p��H�o������N1f̈ҴKe���f��@`<� {�`�|�E�ׁ#d��u�z�i-�^y�Q�VF�������P��73+&�1,jS�S�F��$��Ҹ���Y
9���?�	��
�aĸm���QA������G�cm������4!F�i��@������57j�(����DB6��֩i��Jy% �w�QTpH'��1Nr� HH��)��T �Ǚ�����a��6�vtjg$6�-�T�$!�/>XXj���xz���@���/��ZV��!��n?ֶ���1%��V�<�p[���c5FG�qi^��Q��@��,$	�Ҋ��+���d�y�����_�<gA@����]�[%�?���ڦB!|t	58���L=Nb��-���&d+��6墤���7^�3��\w@$c��rB���"@��$x�'̳�0�^��p�n�?w��)�w�����۶q��,�eq�we'��K1EV�{����(ŕ|�!�VKL��������B����f�SJ�[���ϣ�l���'�3_�r'�f�̜��T��Fw�XF����H6?�u	��*��T;ţȓ��@W~�mN�F��z�(��}�Uo��y�@����1@w���S�y��E��R���t	OYi��g-�4�}Q��� =P����v^&���9r�J�ȁ�&%?�|5'�>'7O���z��7�M�F��G)�:d��*�4�V߱mE�0�^���G�S̴G�����E��6��LxL���C�ܾ�}q�ug���ْ��g#G{u2�ٮ�%�K���[��2~̝G������芺d���P�ٛp4�,']U�<��u�J"�t&�CQ���X8;Ӡ��nr�5�^���R4Sd��������dR�ծ^� ���s,f
���ӽ.�S̋��ŲS4��:��-��-�S 1�o�nn"��h4TQ�qx�}�&Y�{o���
�E��2�[2������.L��ZҴT���"�V����h�F�P���I��:�b�o��q�[�~?�[ą�d�c��k���iCMLiFVE.���8�?P��w�/� 6�:�D�m��R�۸CJ�/�ɸ���S�}�j�D]��FxX�қ8
��I���� 2���D�����x��&�w���KG��F
�*��ԏ��~��	�@�H�!��݈G��o'�p�;&y��&�O�N<K�ri���6DG�&`�>dW7���?�z7�Σv�ɰS���}��LVዏe�7��KR�1�3D�n�X����������_��K�H?P� 嫧���G�(ܩ�Dy��� � o?Jـ��BIH
����LWOK�hz!EC7��$5m�5���ԇP��	m��kJJ���B�T��%x���(e�""EK���j*�Xnӕ�\��$��X��xNay��5~q#,ͅLM(��� ���H���wx�c/��{���(�=�L���<k��2��Dr�r��Kŝ���m��a�=0�b��Z��K��?Iof]x�χ1eS�촙�v�vZ�V&C�&˷��A/�������׊��Z e��g}`����r�����	�X^x�Qc�)i��ˇ�/t���{x�U�f_F��l'�x�[��v:���q���;�����;PǪ��7�6C
�i��nW�G���l X>":��2<���\$��N�����@-	x*(�ȅb�2����h��xƣ��ByƢ7�4���P��h��?�Jb�3$�'������	=M�9c��֩d&��&�>�+�-ز�c�gP��u�t5 �!A�vk��R/���̋��G%72���ǖQ7�:�{���b�?q:���Z��%�+`�`P���x��/��s�3vg��"�����g/�#�я_򹉟c��F�zu9�K~b�?�T�h��������Q��8�����R�D��w����If��2�z��s�"��{���{�݈ddPX� S��]��<���h���+W�*sy�R�\���a�)z����7��޹�,��3?��K_kw�:G�z�����'�2z���ۣ�=bv�2g<�_��@0''�A:aP�w�q�WE�
���-o���d�XK���7�2��i�IYu�#��I�MY�8J+��'�Z*K�eu��57}.[���f�Q4_������	��0X�mN�/��I`!����ON�UK ��Q�YK:���:�Q"��b
��yr�W���W.���%Xȯm�ķ��P�)<��� ���N�8N�<��GP �Tv�3b-D�����k��M���6��4���u�J�T�/���Z��4�1��I_��e�L*��t�vX~W Onm/w�z�f��6LA�q�,/qM�����x���s�[��KE�삎���h�E��<o����o� x�D�D��M��K�� �]��an����R�TKmL�>M�X ��3��CP	�����࿊���01g%WeB�s5�+u�k�`�}���%0U�2�� ���~@c�-L�)�b(D,�s��̥,���{�V�)�ڱ'E�$F,���,#<ŧ=i\���S����L��=���n��!e��`��B�$a更�ȀI��M��W�w8������Iu!9�c��!l��{i-U�c����*+֫ϜRcD�fEpD��PkM�凫��m�}���&N��Lj{��mp|��
�+9]t��3.:�_������ؔ�sk�ܷ�v�����ܿ�����D)T��*��j;���V\��q6$���зTo�K��e�;*�-��WY�~���F�m���|SƗ�<�Oh��q�	tK��-�!3�C
4��J�e��az�c1�gE����U|�0�@\�ׂ��Ǳ"�Q���iQ6����%�5A��h�O~3Jxc��l����S�k�Ck���J+QNī&�C@$����/b�]��M�6�	���Z�`(��#&�͂R�r�lp��� �cH�<R���~X�01-:] ������k�)�{�D�����o�/�w�W3�:����/�i�mllV_���Q��R�nOR��$����'�K�O9u���l�sK�=[��<'�w�oWqdZٽ<#(�Fr �b�������[������l����NԅE�l�J�Ɗ-�Q�+^��^����4��[�oK$rG�`���ls�6z��ϋ���MZ��4��d���@_�`_L�8�(��F��a��s��&N�.r#upADILf������ a7����S���j.5D�0����;l�O"O�+w��o�#<�/�{�(]޸D�ثx.�����`��y7�𒮈���eGk�9���:Gx^�P�)���v��K�������V)(&�>����=� ԃ��ʐ�c���z`|��e�-],�a@u��G��zn7�ݿ�]w�'�bm���X9��1>܃�3�V{}�bJ7O$!WU�c��U2&!�(� 2W��'�V�m���lBB��#��\�����Y��)3����M�������Q�!��D�vȔ�5����^���jO��G�P"gB��	�ꋾ���,��W��m0�2�D��e�]w�u�bI{������&H&�F����=M�pE0�U�Y:=���*vdxw�`�_���ZY�_$��}􉇫�(��M�?�bo�zM�`'�zp��O��ȵy��\�^A#)�	L���L�Yo1��Nb���;�g���w�~:��6���O6��f���j�Ĥ'�u�i�=פ�|�
�/�mX?�A�/���"���Y������}R#�tw���nx�����<a�n����}P���qo��T[������B-����l�L.��0�Gn'kN�TCپ��@�X�Y���A)���_c�Ycr&h5�(���m��@a �P�5��ؖz9����ă"O���Kp g�>y���5�
.p���:� ���|��{�5��˯'���D�_��|�����4��ʱ4�ߩL�Wf��`܉�s���d�.�؀�K�:T���p��ߍH���ȗqfz]j1�K�n5�5��w�کf���L��e���>TȦ��g~:�>���l�ә�.(��M��8�)��͍w��a��M���#�NZv�'���ş)|��D!�º���Im@���h�1D�5���t[2��+T���l�ϯ2�=�+�R���#��{��\@P��� Fq}�f�5��L�8���8�>ʹ����A�ۭ�B]�Zh��I��k�@�X�?;q+H�7�{� l�Km��z����X=�q�E�c�*�N�� "x{���ƄO��3U��Pt�9�
j�eJ�c���Y�S�I��QT�N=�Z�U��u�9���p4q�pX�-�h�~q!aږ.�i�Ηgr'l
*%Na�X81��a�<5���=t���!�{�#|Lm��\�OiR)�Rx�/�=j�&���k��U�$a� ֓�d�O��;���n�Ӥ�Z�F=����Z��֫��:��VF�$��U$�|iT���C(��C;��H��h��$\���č����p,�n�H����12��;����PX|��gl��-Tw����n��'�3�����y��Y��	�tZL�n��H�o��o5pH~�Ƣ@�(��Q�H_��|rԯ�N���E�f��t���S=j���q�e�_�U�]��VW�U��M"����1�'x5��k�J�;�?�GP~�0���~�uD�ꚑ\���\_?D�WV�ū�G1����4d_�3wb��f䜻�K��$�w�^B���}e�����B`k�=��J�{$i�[��	zL��\a��Μ;�t���4,��Hz���6r=�d����I�7��f�1=4{u<$�����)1�>���P �Κ��lz�tFy⇼���Ǎ�g�J�~�rK��׉3��/s�6n�k�P�3���w%�?�N�kӎ�:��z��
���?�.<C֥-�;��,�,VN!�D��B���i�,qJt����<u���֯#�v�PE���� yqE�
�ߗԲ@�-3�zK���Z�	�(4��*�vw0:���,U����q�Qs?V"H�1?2�P5�[�_U�x'�Hde���,�˨H[-AZ1�� ���P[z�lv*O�2��B�2�O���F ��^�-��x:~I��PLH9�	�!���^�o�J^��}��fD�J�
R*�U;���@�TAm�?Z����=���\xe죗���	�l_���qM��A
�/�K��n�RwAZ��pmy$��oQ���Ľ��5�"�-^�]�Ȟ�m��^��M2x?���ƣ3���P:������F��뺪��<VvA��.2c�R�f*p:�����Q\�A��]I���N+�GO�Ь/Q�[�Qb����H��'8dp�f/��J����J�/�����1Myw�z�"p>��OA��V�z0�������q��%����c�����ר��B1�v�`���ήV_w���Cgx�1)/Pr�����ԍ%(�d�?���݄�����*��jB�6���SO`U�w������TpZ�,i��Ṳ"�V`��Q{���F�	�\u%���$����B�x��ʅ�ۈ}�n������ E���^�uVҒov��j�Y�]IZk�	MZ�G��&��?�j�a�ʇh����mxgcY�Yh]g�6.�`:�"�By��H�����6p&��T]}��*����s��b��=���N���54�Ac�$|ۮ]R��)�9����g^�'�+���i\6j���N.6��n�
��ަ�Zj�}���<���l$��޻FI�\d����yQ�&".Zcz�l�ܹEHz5�T�%VķAJ�}%$g����y�� 8E��	�+P��T�$�gӴ"���*1?���`%{�u�!�U�R�ل�MOdb�Qnxl��x�З������c��D/o�s��� �Mk�3�rla�믴 K�ˢ�/�1�>�h�(�Y�d���X��U�����:[s��
@�������T|��0�ݕ�Uٮ݃B#s�o��:�	�7;0c$jLG��B����Zd6? �Ĳ�;�q�C*)�[��y" �v�""'�E�n�a���%}��d��dL��l�=<Ĳ k�����-t3��Ddz2�6��I����*���|����Q!=��u��K��f1F�ъ���)�����h��O�5�������U,����@���m k@;àR�Xd½U�^�}^��pՐd�fK���u�� ������Eu߂ngo���G�Ұb.��a��	�1��OL�Z�^
��N��Gt�p��WO�Ԓ;�ܣn����$��]�tB��J�����U����Hx#���1�D#k8�R�L8�t�-�FY��eиon߂�$th	��2D�~��{٠ pX�ݨ?g����>0�O�`�����'�D��4�����ؓœ�yf�r���j�3�I���dMB/���`���U������򶖂�����]W�lZ�+LB���!V��x9u}[L�:��#�ƨ�.��윯�۹�9x��'#�K�KT�1�<K��z	��������v������҅����"�8���3��Ԝ��l�{��w����Ib����OǢ�b�3��/槻�Dlq&6|ܗ!4Mk!yv���d�=�-t�8��.j�#�k�����↟3kKӫU��?	�4��X60*��Ȇv�p�V���J����}��"�aA6�@c�w�
H|oP�NI��*h��v5�d��/7Ț��B�%�|=����ʶ�Ȱ*8��y����D����SG�|2~��;Ώ��.z7P����1H�X�7�
ݚР����z2��DJX��?H����~'���υ��n�$B%���A5�P� �I�QѴ�͔�U=�=�u�y����9}�ZQ�zo�%]�h��w�'�	U҂uJ���+
#�������^t��ԦUb.�
��[����� T�餮u�Z+�e�b�6]��"����b	N?Y�em�M���H~C�����ۯ%�Qu��<�42%cU������XX��b��W�Z|�����∇��m�<�ݟ�lɰ��u��b���]i/&����D((�<������U�����4�:M���Z��ҽ�P�~�^��zM���<4�A�ض��3:<~�nV$e��4_;�ƢI�4��@@���x�nB�D&���`���������ɢ����1D`�� �k�=䪮^�A��z�N�mi�e"b����B�����OO#!J枎H�QᨢQ�z;O�E�|T��a���Ø�e�'Y�_xO4�c5w>���=�seXbr��j*�Fg��oB�FW�d����;����w��N�(��F�ïG/� �P����IP!�/�O
_?�6-�2!�_��̞��ҡ�0�l_ݗM���n��u+N�ֈ�STn�ԭ{�<�5�c%�M�;�.�[u���uX?lx�H� 3l�����G)��Ƣ��zY��O^�a�č��9<��r��#c��	e"��À��_/����n�8|WH��^��v��h�/�_�q�;[���]f֡��G�+W������J�?/Y@�%	x�Іmf1~ |�;C�4��G@�{u
��C �P�$��"��.�5� f"���ss�B��K�{a���W����X4Ψ��O�G%�Y��Ӳg�^�&O��\�!
�/�<��j4Đ���0��r�		�%%N�Ͻ�(p0�5��6f�*e1���'�%���XV��_�ۗu�R��Ym}#	�z�'�`/L��n���I����H_�l��}�׍�-�����$�����"���7�H1���<f���A%�[�,�z'��h�=Ħ�Y!盬�����f��ٹ$(`�=M�ͲK�:#��(*Ӝ�P7UV{KN9��O�V��H��O ��*=�d+���R
[�:L����-�f�Ľ\��F[��T�Y@GX��:��j�:�xw|�Z��fuՊ� &�hM�"g��]�辽�h!#0 �L��(��!mZ��Ĵ�0�J}��*J�M�e
�0� ޑ�QX��dj���gA��@�|�>�BgEJ��|ch-���p�ld�ws�)�r�	�S~�� 2�|~�5y|sڋV�O1����rH���i�C���[�@Bp�v��V.��(�QFr~x>�Q�;q��'�0��$����e�b�8<gc�S	f�ڀ�Y��|�m��1��Al�q�Ѷ���uD?��Z���|h>��R�O{�/9�g��D�Ey��W�}��p����I�bz���a�Ey�.3�M�f�bB��W7@t�df�$�6�`��Ecf�Xp�T����{=X��-��Hй��7���pHQ�w<L�|���)�)�z��`��c��U>��J �����+���,l����ǵe�<��ٱ��M����X̛�Z�7uXT��M��g.������@�&WT�HكOS�3�ʧ�z���׾��
�jCR�h�m'r��x6�\��E�/�;ҝ�[���xNi�oj�c���Dd@���S�W)b�]Jc�D�F�Ya�Y5\a].`2D)7�)�t`���r�zO0B#\��̵���
V.:��u(������DZ����D�{��u�� �:x�{���K%���"^I����`����B����-�3��^d��W�mDd��R���C����%���c�\��f{+�f-���&�Ke��.�+��h<2k�V�}�M��Z�����z�e�h���&�x��$d4d2<�pZ+h��2�Q�J@�������n��
�1:����݄�FQ9�h���ҧ�Lx�ˬ�I��-؟`&�7<|�Q�l�~���f�����^�U�}*{�l��z�&T�/�;��������V2��1�@n-	4|R�з $}���L|4���j ?�

H�h��z�q�]�1�E�-��e�L�f���(���$�v��W^jnM��+��đ�-΃�S���24�E�H�3����.���s�~�3�uڴ����߲����2;kĮ_K#��	{Iǫ��N��������G�D�_�_�a;!�&��*�SNM6�8���l�nM����5����&C�f���EVk3�-l����3�'�SMT�����D$W(��ִWev)}�[7��<�D��sb�Fy�hC������4p�x�b�m��q�lrG��h���w���ܫ�l�S�xD��R���R����0��Ieoɷ��P�Y.�Dp������&�.������Q�U��\�	��A?�_�t�9H�G����8}2��+���^�vbZnϲ��:��@⚚�H�h�{��oe�4Q����]0H߾c�"�N]�Wr�4\�������BM�^=��숶b~v=P�s~Vհ����{�f����o1I�u�MW��h C��f6�~���$"���pg��͵o�u��q��6҅M��RK�d	�B�T��rA�5Y>k��a0�7d���$Ij�8���,Ĵ~T�M�/`�Q�u׽�掷�����		�����Ѡ��t���d��0�}�,�_u�b^@�a�g	qڳ���8�"J{����� ����<w<�e�'��\�i��2��������5��	~M���y��5Z�".�q�J�g�K���fg����A�����a�P����jGS��eM�6�8����oghm� �Q�;��g�����Mv�k�2�S�Y+Ɠj��3��3�SM��B�6��V�K��(��b߮���7����o37=o����%�l1��k�N@ܞ�u�Y�Kw'�>��^VX���~U&��	�U4Mӄ��U�K���B�ڦ��}��>�}�V	D$��($4���k�Įq
Ud0��ǐdr9�G�RW����	o�=Jq"�\��~y{ġ���+qӑV�	ڗ|T�VR3\�@��S�)P.մ]YK�B`@�
H�o�t�X�#|TN}�����50�1a��`�E�F�4��$8M�2�%�d2?��,Jߠ���u��76�(E��޸r�ԇ���A@�Pq�~/�[���j8�U��x�dO�	Ck���;��b6=�ERkv��#�6$�=3�-"nU���YF��P�!8�[��FLluQ�5C �ƶ�=������tmK��4�ӧv�/�w�Ty����t�k#P[�"�oCY�[�M����Wֳ���_?;G0I22��5�J'�^���Y�Ō����M�U�ʦ�b) S�S:�u��fUࢪ�T�\���>q�|��D�rI����@F�t�>��,��������]M��T� RI�P��o@�:&:}� G ��s�; ��y��'�^�d�҇�4��,�>�HU��-1�����
���Q��}��l����Z�|A��F�~�	?���^�2��&;�W� ��K�U>�˄`� �~�b�&�W�,\2�T���^?�Yj�=}(-�Q����th׌0�;N��A9��^���@�]�א$8�b
�� �!KWj܉��o(��]gZ��؇y��"��g�C5ל�)�}}7W�p���. R�� d<�^����6=�*dbs���X��K���WT"gۘ��eyއE0����J.�e�-��(C���>�S�Y�%�R|/���D�\T	�M �59�َ&��f:噛�������� wMQ9���*U�R��4��6��D�\����N�u��Å�4�L[�S��
�F@���y&�^�ߏ0��6v\�
�����e|#S9�5Z���N��R�|#�Z0��y�~P�^]<�-��s׃�vu��՜�YA�D�>� p��qI-�XY��{��xwV���?�[
9��,�(4�]���Q��wM�U�����Q�2�	%��l�z`P3� ���`o	O!m9��fh������**9P
x�G�u�e��f[����2z�ӈ�!*(�&0�*��F�AӐv��`U�6/A��Y��n�� �-M��zL��xu'���՝�)¨x˞����ڏ-U9�-�eR�zv�RN-LL��B�Z�di�j���oD�OV�S=���o4Slx+=��v<�a%Ǹ�@���D�V|gV�'ʥ�q^z|5�2Tqh�"2q��o�_�x�^�g>)S7"�O'E�D�썌�W�|Z�y������[mp���.'�Hf�(A)��j~)6�[7gM�������+����B��v�/ �p�w��'�5Q���^�%z{h�0ſ&.�[��U�{�}��ӿȃ�R�K��D@Ϡ��Ԏ���ܗm�rO�� )u�L���9}l0!�:ƈ��q�p�ަR��˲2����9�R��iM��==@�yP1�PΕV1�����]��>^�x��ȞR�`�C?���U���}�4X�-w�p}DU$�7A9F�A�y'Y[B��և�l�߅+�բ�a	�Ê��CTbs�����]�\��@0%Jc�V�/�t�6����܎�;k���aIS@�-bRkg�OG�3���j��P:Bڢ�鏇����|��1�g�R�"A��2-�2���y���Q�H�|�p�R�(��s~���W,�AL}�M���l4������(p�+�g���#�Rʘ��l�ި�u��37�-��5��k��xn�d�J�`�(�#|�6���%�T�kfjp�w��®y�k̃?��&v�7��*j'���	kp$���˻	*� I �ȊsW���f��W���t��~�H����!\v!J��:��+�9�D��"�e@Ǹg:�~��#��A��!ϓr&�	R�����T���z�ہ9tAܛ��X�WJ����;14O���n�6�O�(V�Uԕa~�`�q�.XE�Jd"�{zHx�!p �46N���=?l%��9�F
nxL���lg�Q��`{a�4��)�?�C&Y��*�����aE�t´�N�@�F�
�ޣWk���M4h9�t=�PB=�i?�q��SC����uo������������q�! �r� �B��n����*�k���],����u8ߏ��7��凙��ӰM�	>(]'��2^��8Ri�T���Q��D~Z�� �DE1���O�����5J{v��c��oC\�_z�'��n��m����k�,K$��񶿕0k�BY��7+�H39>�G�@*�	��m�l�`�~�k6��.��C47mp���p�}�M��,��*���<X�u��ΰI�E�d�hz���`���(���axl��tW��v�1��kԥ�ϯ������[�^��`�<��*����s�t����똩=C�ßX(�JP���n��^�ʙ
���z+�_���h�^���0���fv�\��/��G��ے�Y�1@_��Q>�k�
�|U�Rz�E:����u���IbD���f�R��<h9=�q��z@�v�?p=W_Sp���9EQ �,��|��w
��O���v�o~,8�A� _�/֤@��Px���v<�T]݃��Xk�3��S�3���u��N� �2�#v`//����d|1�� ��m����#e�0!]��x�#�0"4=^�x�]k�ȷD��೻��@�o524�M��6R�V��^L$0�����,�e�f��.���X��G�z:���<ڌ:���H贼��GK`�O�3�����{1�y��a�w�-��g�T��v�A.F��Ǝ��g�Wc)�B��l��|]\���I����� c��^=���Л�T��:�����-	�$ ��9UB��E@i�h��~�<؍�I�h��߽g)���`9�["P��b�A�^� s�1��!�6!����-䄌��$d���D8y�f"[8%ģn(7��~� ������������:|�c_'PXcP4�����mk��]외ƭ��m�����Y}D�<=��|ͯо(�z����-ǝ޽0������E6]1���@�hK*��#Z�-��Ϋ_��s�k����bh�U���½!��A�Z�,7g� �Q�|�JPtaL����#8� ���P��õ��z�z=����_�Z��H $n]�n@�1Pl<�hLI[���l��U(�w���)3D?�����g��c0T����q~�L;�Kp�������A	-��AjLYg79���/{`�������ؿ��S�e�0��8�
kh�w �_ ;���K��y%�\e���✚^"庝�U=6��Í'�����ұ7�D�R����Vg��@V8�^U��Hu�B�6�\�?G�Ria
�N��)ND5u�4!=�d�8_p��хN5����9}�ZlHP*��w�45�s���0WR4�L�ʴ��Y�<���1��_�3�����!�<�6�+�K�������r�b��W�i�cNj��tsXg�+%������*ѫ���&�b��	��;�;���$�ks����q��q]y����,h-��l����
��,��Gg����`n������H��j�_L%���__˯��R����U�+ͰD���	�v �H�ž��6�9ѫ�Κ�H��"zUc`�W������W�hѵ4��Ԝ��M��7r�:��/j�ʬ��0<,��;�����OŹF�WK�hDn�P7@�����X��I��0���H6�XXc��c߳��}�9$|���(w���Y�GU;Bd.����%���Nz�oa4�� �)3v��(�+?�����h�9ea�����{�{܈�Y� }'唠*��i|Rw�Í~<C��Ye��	Y`ÿ�r
���&ڍ@���/�"�Z%��՝�5�"˖����=7D׆�M�h�-#�������ũ���=&!�m����V��G����(W��6�K���go��a�.��q��ijLct,!R&m?6Ֆ�o[����5��B
�~ҏ��Y]�3�wO��{9{x:��	����vl豩��C�(4�U0!  ey�D�H����.����W��������`�q�Hj����%=�!�#n�G��u��N%_�r۳��(������S�����Lƀ�eS�[ޤ��H�APŎ;���E�����D�5���A7fPRD�L�%ɽ�I\YqW�ܸ֏�5�v�8w�]ǚ��a|t)���蔺.=���v٘�(��O��μ��L1�"����*�Dv��˔���Ͽ9NN�=�v�f���������C��pc�X�PL>��*�[|� �9(3}3�	*�w�%�W�#qx�K:hٳ���Uh*pT�?^�%��C`5(��D'��8J�6�T� V�GK���= %8d@����O~ziC�Z�g^�I1�9�ڠ�vRQ��Sf<e^z�H���;q<���}$��uǰ�l�Z~�Q\�����U��
��yf,�A<�K��~
�=Z�B}:N�����U{�RW(�u�q߯u��U��5Gi�s�OZlE���ȐS�d��!!܅/U�wj"�U���s\��0.�8��f��YOn�ݭx��V�?�ZwK8(Ї���=Gk�J��s���B��.� �._��wx���D����� 5p�,s_�1���ˋ���@��.�R	p2,�*�\�^�+�B��k�K���A��\'�H&�"�a���T���+C��NcO.�X ��a���`̅�݀ש_Y���2X����<A��l��DYq���X����X�RO��B�i��d�'�?u�`�`9F��%�����ʇ� �B�w[�Ր�YE���yZ�Ki��T� �Y��~0��d�D��b��
�9�Vt�/YQ(����%�C_`�D�gr����}̄0�;���Myq�k�q��y*�"$���O'ik1�Jjs���ro�0~�tѝ>��L��'�W)���#�RG)��U�9�+Yis@��ű��#���iz%��`�����Q�0����{)@�q���~ט���LD�O�s�K}�	���M�K�7�5klE��&����� �=P��9�l�UY�Q���:(�Μi�:��,K~q{Hq�ND6��*�a��%�����I���[�gFJr)֊���?����L/(,���u2�so�4����.;P4hӥa'��5�%O��`� �9�ς�e�:m1�qF}3�1���곩P����`�!�� ��<mC��N�ѳe5�U*�Z�H��Q��u��-{��3E7}GJ���	���?L��f  �W�
������B��⚈�M�e�	���七�'�\�!�"U����b��2��̸2�ە��u�n���.T�N�23*��ЯC��?��l�^�N
�8�nz���K�E��a7]R+<��%]�x�s��لߙ�9���׵��rS��q��3^tB\Ĥ+t�2w�J7Y,��q��6~��L���,��������R[�#���?�Q(��+�v��|�B��v������jt5��}���`�h���O �;FGJ��S�����Z�@��k!4B��bY�Ϛ#p��>�>e��6�L[��$���Hg?+W�xƆэ�j�ޔ����x( (��⧇�������1�gUT�&���N�/�V�^T#�i�.\��Q��D���_e�O�?�^6P	�b9�d����{` M��w٣���>F���~�O�tq8j�81��)�O
h�l��f}Va:�q��3}�x�Q�60OD�tEu7���6���p�X��s�z��P�������k���`Zx�R�
�+�kDf*�,��C��b))F���Eȩ���0��{��xp�l3۳�`K0���p^]�мd�~Mڞ�鴊�����j�6h�r;���q�t���5�W��IY�}BdS}�HiR�(zn��4T��=e��D�e��ME�=`�P�"�!�N�2	nE�V{+g��<����͠м~f�8K��7T���������2ז�	���Ӊ���2}��YGWb�a\�A[S����>;pw�0�x�V}Rg߹
�����
$z�V�k���F����� ?�	1��8�N�..%���K{?�8zq�1`��uLJi�⪝���l��)*Gmo�_y[^^�)�B���G�ih�%c�����(���?]��i@�Ũ
�%���Bv�;0�%����,�§��l��2K�4Dz�6����ޑ�E�ǚ���A��i�/���QD�k��7� ?0Ā-���TH�����=d�sv���kا�lLxq�E�WJdU��*cuф�1�Pӟ���D8�]��H�R�E����6~��x�����,�^66
)���@�h�M;�$ �U[�B�q@@�=mb�hłS̳�$�xG�UO��XfHS��?F�|�'.�U`3���`���C/Ea���7:��}��ɺூMu8>�s6]�G�N��W����z!7.z�bZ]p��}��.�8�AU�٫Y������\qY�<�Y�1��Z���T��{�֊8�S�p=���Z�.9�������@"f�ζk�a��o��4�K�(�v۴��A���c�4k��L�:�������^kD��7{�S&̵NE�鮀��%�l��[��N�u�E�b*:k҆U���p*J���W���Զ��lm
?q���	�G,�N��nK��������8�\��'FY�3�y*�=�[��1�Nz�#��<R�x�E��D,UC�ڪQLj)�7�91-��DG{�.�[U�d�)]#맨��TB��#O"�������߭ڀ]R�d}���ƣ
���?�+���m�lSe�d!�b����2;��_� G�.�[~H1#�	��q�N�V���0�~�5�"��rJHf����E��ΑAH"Ԡ�3Ó�Ra��Z]�"W3��p~�t{`sD���f�_���mn�,���L����6�.�bR�I��� ��Zf$�B28	8��:�
�?�n��R�DK�ca�����*bͩ<x1��,� ��Vh��T.�7�Fd*Ԇ�.��$�R�&�0��Ų�����cB81� Y�؍P�N�OJ:еi�u��^����^ш"˗�H�lE�WZe5��̬�˼��5��4.�$܎]�
�؃�Ǹ���ͼMU��],��[�wJ�2�.�RNLydfP�͵���C�M�A5C�J�]O蕾0`��I3";���byw��]�s�ݽ.��)�#JC?")�.<\��l2i�e.���5�Ο�\̀��4�',��K��� �B�<�>��R�(j�.�=鑞�-Og����$c#���F��o۹t4�Hu��̶�jG<_��y���>6�M���/���������iBR�SsmF9]^<4#�̞�F��L�z=�)kT�5m��eK�(G�d��p#~����"��%�I�kEa0��t�P6zHߴ;�'���m��J�č�@�	yT{���1���	v�Mk*���0 @��m�}���PNB��7/o�bM.-��@,���h�ć�,�;�ߏ�%��CqoQhTWv�6s��Y��4x��$]���q�e�lF�&|�Z��h����`�#J�'�4^��sg(�8��<O!�,0s0=�|V�\.(t��Pt�ǄleK3�V,@�mũ��<�s�|��@��:*uG���߅I�ۈ��Z�#u�	����A��S�I�b�Mś<��+�@]�ց�W���~���� c%����ĎyeH�M����] ��n��0�T�7�A�oW����g�;�D���Q�	�m~�$�X<���vbg�/c�N3Ē���\0p�pV�R�Ae�8�X��E߇�i�xg�QGv�"t׹�ξ���"�.�6m���+n�&8E��.,_��H��uF�����	���=����R�!2��	y��v��V�߲�ojp��މ�"�,<��3��CE�wc|D�5�g�H)E�<E���d4�^����\3Y�ZY�8�A���%�!j�-ǟ�h$)C�Ps��K[ɺ �]@y��aTB��p�z`�|J�՗�Z��W�1Ԇ�W��t>�k-XP�^��p��@����>��f�oa��&m>#Ě�,/�*�m�сr��˝�ʩ�����AfM�گ�>s|:!�n��q�f��R/3Mq08�ou�"�=n ݳĳ������V�o�R����o����jT�4��Bb�O~?�T3g�p�D7��f�������f���ϣC�
����Q���@��6b1$J����ל���SLc�/�}f��K���v��;�����4D�����W�̲ڳ4�z�,�D6iM��8�t=��y_d22rb���G���X�ʔi�����b_����:T�:-�f���ʅn,Y��鵯�L38_��b�&f]�+���覷�5����:M�'G�e�E%k|+Hau�Lt���s�ǹ�I<�S����MZ��=J�"�0�?�QθO'�3^�n�E-�`G�ͮT�BO)�V��Nu����m�ʻ�G�pi\ ��lh�9~�קĝ^��:S蝷��
��-Z}�ӫ\$�P�a�7�����[m tnMOZ#�WSr"!���5��%��Ѽ}�uF�c���/��G�܋��8�ޑ��k��V�
R:Pm+���,�chg�����K�ʷ�::����qC#���f:���(qK7GY������0�yߵ����Lc�˺����d!z�0u9����{������C.�*sq����6hv0Aޑ����l�b��z�}�h�8Վ���峸��ntX��%�u��C�\ە.P�*�����TQ��rA�B��q@yO�2I����!Z�������Ȋ���6x��7����rD'���4�����u�{t!Ӳ�pz�����Y��+����e�:���3Ie�$�<��b���Sg2�v'���D��y����Z���@HT*._?M[;fO����@���2dJ�ե��{{�R��V�ZP�X���
�6�|.̢-J�i�#2�dm?��>Y{�$]�V�!����L�<|�(i��n,�>X�m^Q;�n�6����e����>��Q/����&d�����e;��'-
`0?L�ߑe�X �_s]!�a�ڼ�8p�U8��ݨ�pλ�CE*�l��f��i��,�Μf�U�<��5V&G����F����&u��-S:�d(��77R�aB$5sc��$�GgMz��.�Yz�2ǃ"��I,���H�_F��}��i*^�H�9��Yn5ۣL�u�adfB/�|�'ux��v#���wأ��Bj�k��`�ڨ���c?P) ����m��2C8W�Ty�.�J�BS�*�ar$|�H�z�?�U�ЫJ.1� F�ج��:/��3
���X�d�$�%��u(R= ��i�� ���K?b\y<S��(�J����*�"">�o[Ap��p�)ܶV��!�+�	�?!���G���L�Z�W1s�ê4x��h�Z�UBm���{���֡��NR�C�ݙ\�)kh���!A��ik�-�J`�
^7b�%����N�H����GR��s@Wa�kS����&�x�#�:��j�K�=:z�$�����$�^��Ċ)#����1W��H��Jo��]�qB)D0ݙ͒���cw]�^7��e�"m�(я���<���1D�䀰�6{?�-Y�x'�!Rh�`��bl9l�-�.��&�]<*�]B�*���Tt��s����Q�'�p-ةEA������i�*^����Q�_�kJh��-��x%%&���t��g�(k.����2�-�xs`���UPH�	���;t5�
��|��o$	-3ZY�[� �TNJ~--D[h���f,i7��j}.Jm�K�Hl��$.���*-�<6"�|Il��jɱ =�s���)�F�x�!?x�8��'"�z��jWf� 휷�L�(%9��ہ�Մ� F�֏��"�֡sY:s�"x�8bhi�u��ܥ;�nWʘmr����mS��*���rZ�Ń/�#�K4�bŦr[��
FǞ���ts}��	��@��������������N�܎����Ta4�OИ�L:�1��_epD��\p�q��m�� �GIXǡ�;�=@}��R�Vze$굈_=� \aa��|���Ƿ"R�;����%�kVo98������&����x�1�|�8g[����'%|�*N��neĐ[���$��g-�����w�!�0��qW
rP���mT��`=o����`�X�>�7͒���9H��M`�_�Z�L�W�U��^cd��]���v=����뵓�zO1�J�P@Í�P�2��������BZ�_[!家uwpsW�>��mU�<:�p����*,���$�Ca�|y��)0[��Ɩ����o������y"�=e��J����T�L�W�x\Vv�fE1��[6��g�Pu��[Z�����7⽩�v��E��o �B�l7ߛ��$�i�=%�/1m(����[�ު4��Kd����d����L�^+�E[QW�� �;@u���S��d�aՍ�Jgt��[8]q��:�@�`m"R�}�m��MN��"iO������E�6��{!��) ��(F��F�:�+�5��Q� 2w����dr�3rY���� x{��$���봹�|�
Į�!QK\fx�Ʋ0lS�)ꎐ�x���"�e]��J�y�ظ�'[8���\�3�nu�em{6B����"�R�i�b�������=Y9�R��B��g���~���j^�|T�Y*�< W���-1(2 P�F���hF�Kh*�B9����'��M��l2-h߈����&Ө�9)�I����	���%�tZO�<#�.]ME&���TH{ir�v���7[l N()����8t�	�K^���1?�F��(�h8�K��I���2�LF,�iB���j��X�洲�sY���{0���	
j��>��]�t%S��n�7u-Gm���O�%���ͣx��rmF��a7?X�k�i$�7���A)��t�$��a���R6�恇ȗ��Uj��9��j�������-}�M��i�%���e���3�J�&Ĩ\wEO�ߩ,r��(6��	יn*�^�w?[���tR?2L��J�,)V{j�82�Ѯ�����7�!�Zj�\�E\t�lbma�w11bM`�bJZyޜ� ��1�{�;�h�Р<��G�a�ؖ����Gs8�o�5�tcЪ�y>Z����O~�i¯$y�~�v�W��z�p�S�";��9Ng�?k�H�JWn)��_�ۀ�������i#[f�=Up:o
Fq"���&wT���P�fJp�I�'ս���I���7QP;�$�f�pw_Ӑ�{9�PM��/8:$���Ȑ}:{L�^�X�P��������9�߻��ix�l/�I��Z9�5��
	X����Z"xeг�+�ڥ��9�2��C�z�n�>Eͳ�*]o�+'*ꤜ
�\+�D��I��"�r��'&]{�c�@-�Ni�U�:;�P�8�L&���r8����%n���@\����[J*6�YQ+��c��g�X��W~K$kT�
Z>���������ـV�{�U9�7��&��n3����B��о�޽Ut|��1S(۶�/����J2������u`a�u<������
�3�I:qٖ�;�ס��I=��jlΟ���bLG�P�Q@�[�1��w���_8[�+ud:�yBrb+�H�L��O���*v��NN��(��W���� h��,I)8-3�"��П�H���#w��WJul�}���v�&"t9kЃ��D���{N3+0�K[�e_��LT�+c��v��O�h�I�����M�
��w�ԏ����T|���<�M�������e�.��=�ʧIί���]�����֟���p��Bc��I���>��w�;���t3�p&.{p�����[.[���D�mU�l�w�N�s���F�2^��*s�����|����	mO�kMx�$���+��N�i��+"����`5ũQ�e�7[x�t��%��1!=��Dad��m�[�������z\_���Em�����U��eQ�p�R�}�0-t`�w:@e/>�hE�u�"�k-�;jr��?F���	R��ơz�<�S]s�l^��Ų���|K2��z���ّ��9@jI�x�2pS7���G�c�E0|n]4��䨭�C�"J����vyd���|Fm�����R9��
ᕇ3h}���|�Fu�1/ۻ�	P�%��taA���1Z�%�)�t�η�s0wm3@��}k=¿��kMx?ºtP�2]�����0�z�_}��u Uo��3k�o[�EL�mw��|���1]^�}���u�E�1@h[F�����hkU�f����G"�6N�.�չ0 ����4�1&'�OJÿW���1�=��(%�ؼ�t��r�[R-��}�׾��a�0���SP���0v}8}��!3�x�[���MFC1K��//�D�������f5��3��7 �W�0ҥgἪ[-X��P{�<ۭ���i^�'S��Iz��'�04{%E>�Q�8�?e��B�|wK>����׎9:�o��E(�XN5���Av_� 3m��]x�������\��,��\��ǀ@_�=0꣯,0�{�0�/~h���T�p���Q3K
,`�����(Y���]S�	m��(: N��8#[\�P��*#pާ�����F?����;��������k����f�fY�@�dY�Kv����j�6�K�Q�R6��_�L�+J�,%m���;fa��EƹMK�"N��Q��u�!��R�]����)]D۴��w�$XB�����$)>�7������~��
�EQz�/��7�|h3��]�ɾN��5�T4̾mP��ؚ��q{V���i��4��0c�X�	�O/�����S����ε�?��F ��"���o��q�PY��@[y��%�������v��������Y��Ёu/TƖ�Y��E|��|�!�b;"�V�Wg�LCS��7��]с�^wb.|Q����d�[HB�Î݀,��� y��	4Yחwl	O� k:��7������ժ>m]LéӬ`F�S�k����JM��إ���j ]�B\���C.JyNK
��sF����(5��ᾜ��`��y6$L_�3m����㮺 -�����l��b��V��W��'�d/�F,�8S'A^�Cs���-
�hx��.T{/vʍ�Y��t�t�Rռ��L�01��Z�8g�`u��>>ig��R�R��p�2%���8�Z-���Aq_Hx @aD��	�tX�o1M�\�$i��cZ�|� O�koK�S���i�-`�E�|���U�4]s�E�n��1�8�����(����Fv���4s�8e?�r*����''o�m]g�-,,�Km�&e<��=j~�kz���5����R7�4�`:����@v)�X��4L89-@a:3�'��K^'6�Ԣ!{3&�����t����k������Ĳj�p��N�PJS[�w;�F��|�:O��w����<���suJ6�m����l��W�x���	$uC2����o��j�U%��n���; �C0CH(��:��Te1 Ճ�l�ܖb������#Dp� �q#���Y�sZM^&��];��:<[ݴ�8&%�ĥ�(%�"�iKr�ש�Y6�;�}�,ѕ{�I����"�n}i�db�E��(��2��Sz" nٽ�ʣ�S�$]]dc�tɐf\��}�i�!��v�-�^Su*�M@��1\<���$nۛ�n,u�XL#)�fg���x+,}h		��}\gSS\l�.�9� >�lv�����5������49��)JL��!�e'/�٢މ�Ex.�4�z���4�0��|��F'������I� ���@]�;��aH�m�E<�!��_K)��X��2Ě�7����!�N�9��
��͌O2l�d��RwOl%��\Ps	(	��y�"v��u����
l���`��>�cH:�:���4^��v��M�XM�|��j�߿o��(�F���9��:X��*qT;M+��N)ݧߴK��G�I��&��H�޸��#�65�d�T�xM$����BzZ��m3љ�aڅ����O�o 9��aD� ^��CܫF;9o���:��7��u������.8���"M=�o�-����>M�#�a_���]~i�m�J%�%��g��Y�6/�h�,wzr֍н��½�>�]F$i����Ϊ���8F�ǋ5Q��^
��ՇE��S�yR�ZF��w:XnA8����gx ��Z�ekR9����U�! *�d�9�G�xQE�WD���E"���_e�j��m24kώ�zYu��q���H	���̈́*Ć�T�FhrxiQ�Ç��/R�SLj
O7@P�ʄ3�.�%1EĝB��@B\��#��`v��o8���ռ^����E��e��j�*�Ga�8hoڍP�=)D��3��Q��b������XYNo���(���Rrl9魰��������x�J	B��p���`�/���Ӓ�Nl.�]��83]�Gd�_����v[c�<�Q�����X�'~�,=`V[�L�^��ß
�;���n���(Km��+�G?_�&[܄0J��K��9�X��-�]?���¼�:������z�+V���:3�'%d�@,#}�m��Ѵ�(��Q��/X�fQ�Ո3�Mu��DsN#1��$����Xv���b�T����P��-�kX!�]��L�L��&���ګ��49� z|��Ms0}]c-K�ݚ%��Z��Mpf7L8qa�����Ia�L��3X��È�{E�d�2�1��S�W�p.��?���s�j��1�H���F��vh�<�^W��vd(!M��B��t�>��9(ez۔��V�K�2d�Y1�E8�f���,E��/�|�@m�V�B�����i����s#V|5"B��g�?f�:������A�2��nJo���
���'�����r�����sG�Zk'�X�dq\*G.��#S�]r�jHj0��4��������Sv-eJW:0�P!y�[P�վ�{66����I��>?��,��j�js��H?��$�O!o�x��׈v������QǾ�!j�z���6w ���\f콕@����~3�
!��X�K�eL�/E��-M�+.x����
V+���c̆�3��pRDrB��a'�d)�k����e��mۆ��n":�.гےTe/�,�R[�)	��޵a�y�,BK���U$�m�z~�����%��v`�sSt�_�|7�5�p�b�S�C2T���������&O��\�HD-�(bl�vXۺW�յ����#���dTS�����kB�o2�'Y���J����φ��o��·e}��EN���&����`�n)e(�蹆���tW�_��GFK�1�m	&��˟�u��92Ӎ��rg�d�p��,䘟��a�E�0		���ݧ;"�W��߉ܱ+�\�X��A���i�����ͤ�G�p�� J�sO�����6t��D����ꟍo�>ih�������t���S���H��@�Q!ˢSR¹���
����[#�q�iVdǺ#r2�wW��e�F��@���|׫M���,��H�I+�ܖ���z~jq���R+Z���A䊥�>,�U����i70P�=nh �����Z~��!�q���F{���G��#	��K-�6�3���@��֭_[=YB��~b9ÒU�пL�p�Z�%�Ed�MP3RL�)�r��k���c?�� 8j��=I�v��#M�
M*4���Q&�A!��W��� ��tu��	�m���&�9��$Pn@?v-؃=�������|M0>W=^ä!ʗ̆u���)9ԩҫv�Ĺ���ד2"�c&����`[U�g/��lƭXX�ѱT�uN �	\���a.ٴ ��RM��� �� �r��t���8u�����v��QY�ۘvL��4 �l���Q}�j�W%X���2ߋ�,�}�W^�B�/��G��[o�I��8��A�h�6�	�����`���|�Dʔp�}���(w�m���E�͆�=��<6+��䆎�{d�����11���7^4�!�v�<s�fu��TS�z�嗅������"(QAT9���^Kg�'�� 0�s^z��B�>��!1�䰪3���$~&�Ѷ����T����O?Sg{6K��xd}��a"�ù��C�j���kG��蘒����.k�m��P����V����C싩� �6�t�o�Y����Ǔ�DN2�c�`z:5RgB'��R����;�5���i����"�{���4���<s��͘+�?�󍷛��u�nGb�Vh'X�	��L�Wb!.niF�劁õːY�b�[���^?*���E��`� W�����LT�Le��t�����_��w�BpG�=I�j*H;��L�;:�� G'�^�\���x��.C�{uG��FFJ:WŪ�.
G�HN�|<վw@M%W]s>�g�)<�m�[~M��D�I3��uSWG���Q�c����;�+zD�J���\����l��9�5}�����C'���=��P�	bx\�B��JS�Jg;n��Iw���ޛv�~2�O�h��MW�f�<�4n".�1���ȿ�B��ϸ���r��O�sR�J�d��J7��7R�O~�YH��F�n@.v`f�Ҿ��]���L����	#laD�`Z=p2�Aed9R�3[��N�J�>�����,!�`o��a�y翧ޫM̨8����^dG�f��l�3b�I[��G�Ō��qo���lz9��,ṛT���W�5Zfr�U$�j��|�/p���
�\�x+lg��^�]k�� B&[�,.[K@��E�D���IF�]�Y�O��d�q�
B�cr#:���V�b�		�G�STWn��t3{$+�@��)���)8:��~q�~px�x}�նӰŝ5���Rux>���0�@U�\H�<��,&�:����Z|��Ys�}�o����ѻ"��Z�8����2cc@��̈́aK~�!�lz��]��<Dﳼ��C�<y���^�E�f$_�h������0!w�y9-�r�-�|�V��\�d�������d�E�\��*�{� ��)_(n'=�n���^H���[j)[�A�U��z���rӯ�j��f<�V��f5Kt�U������-E��l,�K6�i7�vˑ��+O�U|��4�''o���kۀ� n�t)���7�F�-=�k!��NI�2]��8�;s�� �u��P� �����yn�R��ϲ�����by��b��-�(�C�at!Ci'�cp&V�-����۰�����gO�]�O����Sƿ�j��rw|w*'�i��YV7��䈔=j'Ǣ�OAW��#\��wAX�]��0����(0j���U��ņ[�k�-��r���Ў�6 �L��ލI�7֤B�VuV �	���4k\SbyM �������~l����������Ot�(P�8�ތsp�Y\o��,��oV=D�6Ub/�<}�������^Ci����S��ŧ;:}4pt^��4c��K\h���fs��^�_��A�7Z*b$�"�a(}\8�9�����N��4��VyP��d���$�f8��L���������x��L�=�I�jI�>:�m3ն��4�[ɒt�<V����8�p���$�HB'/��#j�A�"@��I���!\��]���D ���)Cs��s'X @��n;,|��F6��HCcP	�Ϋ����������G�BE�����@�yVhYmC8aux��I�"�Ǯ�3�PC�7r��9�іt�����k^��v�e��Ɲ;!g�L�L�o}pb�����Od"j��?.L�����V�<N��X���}���/�*U�����ch¢=D��Wj$^е���B1!Q�NEٯ{xo��s�0���<���D�:�g���N/c�%���V�hɡE�4�3�-̦���4�v�߽&qٷ���!��]	"��o"e�e�`��T�a�?,N����J��^}��w�s�@x�a��׻?�-�X��Q=]��z�`Y�`�vi���~�[)�٤v�r1Ý�;:��E�gsv���Y|<�T"�y�sD�kΎj.� �JSW-oA��? ��k�O�h�Q�ͬ,X�N�8��1�ѵ_~U�!��|0ەV���Ѐ5���2 p���֧V�f��W�#o~E���f�.	b!��	�0�� ��{4����O�\c��3��M[�ש^*�D�2���d#����tI�Zư���K5f�篫�
V���_m���^Q!���S.P���
����A
��#b��M�⧐7Fi��<�.��_7�������4\R��?8F-�l�>Py��deE�o�u�(��x��G}�R�ڄ��ޠ�ϡ��W��z��t$^i�Y����d����OiQ�%�����*Z 6`2�k����#g�mq��WmZ�PL�h,���m�$̿<�|&X��~�0��t	�y�sQu�J�}ۡ_$�'�jV7�+QQ�)�hRg
 �d���PCz�(������6.`�O��۴1�8��s(�H�1��Dh}/	t�*�M]�e� #�F�`�]���f�(ݪ������iT��k��B��p�c`�dQ����<zb|;�N50��	p���6�S��i*^y4�i�C�HR�}�i݅f����8+�sE���Cb��2��w���z�z���}�C�f��w��\���������5]��(�J��4v�[�B�=2B��w���K鉡q1U�;_�ג)?9��w���2'F��,����p}�����������t�~����nw`qY��q:�h�쯮�z�9�
"�E�
~�5<e��i��4_W��3���/ɋ�1ek��X�����<lVs��P,�������XO����*�b3Cb�z��뭱B�dvK�3��$�p���}}�Q��#Sw���q����qg=�!�M�l�'���~o���Ԧ�E�0=U��!O_*PK�b:Of�3`u��lf�"Kc�J��&��u�����q*HZF��%�Xm`�S5e�f��M���ox�X�C�!�(�-bp?a�a��`]{��ޙ)1_n�rh��\��]�_d�Dh�̴b ~îUZs�n�Y���/U�Ѹ}��4aO]oj@��|3��>�7�qQ\�Pl��&�uveFټl7�vO����cl��H��~��^�m�%<���~[�J���dD��3_^����%�BtG`� ��b�%ry�jӟ��u(�`�Q.Q�����%�s2gSψV6l質���҇CX��ƫ蘡-�vc:�2w�p�hi�n^�L�u��M�����Pv�H������ybf�����j[�������=��$�J�`i6���8�W}ug�6�� =�&6�a&Xڭ���*3n���鮧å��ŷ�g� 0)���k]zڞsSi��p�<`�i6�~xY�OD%[$ѥ�d��8|y�k����iZ�C��\�}%���E<���w .�MRv F�6�fyP���Sak-G2�����I��ڱ�Ko��/W�B�Z�,���H���~Z��zwW�*�q�H?�n��|	�8苿�Hd�.�p��A 8~�2�����C���]��f��/3^Y��3�3X)eAzu {��K�5
B��o�3	^ݗ5��iu�_Ic����-e7fZ�:,e��![(x_5r_�	H�[�, �P)�z#@�Z�L}���3���
�v;����F�x�s ��9
jwlF&���o�OΙ���U�Ȕ�8Y���U�D����o�nT~�e��V�ڄ�W,��<Y�$�FB#|)�RXL��=L!n��+I(�%#o���Xm�6�z�v^Y�X���ASkir,��-{@&n�&V���o�P�7.hAS}^h^`���l�N$G�6�q�z�Ǧ9�2r�L-?�>e�rN~��Q�i�I�(�����>5�8�\�.ؗjD$L�[�Bsb�D�Wpz�����g;�U�j�ΣHrXp�<\��_��JT�)���x���OT��Lk=h� �j%��lk!�Tz1�M�A�� ����NM�Z��D��,v"����n-�zV'�m��1K�`#�b�o���v	�j����Yxٳ��"sl����r�֌3AIٙ��Wc��ՍP�}�5o�_:�lݱHW���04�RK��ht`���y����
�iL?�E�<�2�	�������L#js[b�P��˵���s$�һ����8�/A�\ft}����|?weZ�����\��Q��^�e���Y�[���
:..�Ϟ���v\�.R�<�wI�hza+���QrZkr��6 \4pҔ�ef�d�e:iv�6B�ݒ�d�lX�Cp
�M%��1�i���v�@т�Q��	B	��#Y���W���k4_u�nL>w�z,�����K�u�
��g�1��%p�$1����^�t�>�KƚI�O6SΊX���'��8
_�+���3ʌY��������ЋZ�!*<��{���<-��]	�PhU���4YS$��h��Gû���.�$ES�FEv�#d�,�n�F�Jn;�\���#���{�dA0/����������= �̀Vɤ`��.�TY���]� xʵQ�2?Z֎NX{�r�]q��Y~D�7�)Q���\-*�m�<Pϛ�d�2��nPD3ZX�)~:�� ��(Qs6d�$^��v���_N\����ڦޏ�������}�2�}_8�K]`iyUds��)C�w���܍�m]����[[�;�fe�;��F�m�ˇ�I�S-�J�P�����9�xxz[������Ep@��@e-��L��1Àya���_Mj�������2��x���)�{�D���-��Mkdd��+�1�`�u�{E�@PQ����<��d��Ƀ���{��*�g}l���W���}A��I�Op?���n�c��y<Ġ���@��<x��8�O�f5���I�����V$X_�U�O�e��E��B.�=���_�m���¹��?�.�U��TR���%�dLg�u�H�]�`�/6)s,j�{4c3�����|�{�ݬ����I\e^.Ml��JI`�4�`
M����m�Ό&f�0v��l�'����Ya|w��;~��w1"���%C{Ta`��?<,�����W�yJ�p�)��Uȝ�8�Np����ɮ9��p1�:>N�#�����>�x���CL��3�ǈU��H�_%{�8,�(���B�à�QJ��j���d���̂�gMA���Ӊ-��)G��on!e�StS�^��̥���~��(��݅�v���f�QIifH}}j�|��9�tuU�T��p��|�Y��K�vA�� ��q�r��W/
�mN �l�K����V�Wp(q	'�rp�RZߛZ4
��F��������4�%�j�S��z�$���EկR�k�Z��Pb�9F:��j��(ަ��8���
�}A0�}C�{��R���d��x�<[�����<[�G5Ʀ�:Y���K�8��M�W�_���5��M5�w�ȟ��{/b��^7����p����(��^P�������\�k��0��E֛y�Jy���<(�ź�Q;"�����9k
i��X�V\̞��&"�L@�0&��X cZ����џ�(w����JTn���ag�;2J"QH��l�8�D,:�_����fn��y�'xܼ9��ȑ��N����]z\����Z�y7C�0w>3�"O�P�w�X$b�/�1-m �Oi��<�)�=��Hw2U�h��X��^ 	�nS��\�)%������ ���[�%�08�C�Ų���v�w��-��!�p���Wc`�:�i�BOh��ɟxґ+k��Ǔ��R�&b;�Y��o"�c��d�R��8Gok���������c> N�o$]g���l���Xp�h��|eW/��~�pޞHKi
��b�
Vгf��j�nJm�d�7�!��"| ���,�7�s)@������,��Bnː���7~|@VU��*�F*�Ϲu�\����B��E'J��P^:��z204Ó��7-Œ���$.6�f�a:h�DB�n����˅Y���'l�f9k���1}i�ur���t4�{�CK�;h����2�=i�(2�SGϤ-�EVCtB�H_.�S;����΂^� ���D�>�c��ň��D�DK����í�Uޑ��/*n��DB�/µ�Q���8�R�sA���X	��®=���:�=�aRD�睷j�[]ρ���H:��w����1�l�?�m0%�F_5ʁ�֌��3��j�Q��0w �k�@��H
	~b�+�pO;�D.�m��@Ѯ�3�+v��^@a9�Y{6d��!]o���Ɋ{x�ȲFM�%V�����d�N��Sg����"�-M�t�3ҟ���Y𙱴щ�%j�Q�6��8LĞ�|��/Hh����Hg���&Բ�=��CQ?�����Z�â��5ʌ��E��o�,��"^�O�
KJa��i�ۛ��S)i�� �T#�3<����?�Q��H��}3���W`�O��"�����f,��P�"��H�gq���=����1�����Ce;l?k�d-��I(�n%M�������Ԋ|/��2�O�<��B�;;�����G�X�wN��˟k'`�9l�P�$�[��;�[]%�԰�b[�������Ѣ=!/M��qI��1O�*y�y�ʸ�}Zy賗�{\z�`I�W���Յ���@uY_������7H񚔉A?�?�+4L�@��,/��-�痾'&
YZh��uh(��H�l���]p�uTA�8��	%���e&~3�N�US��@1`���,aC0����j���E�.E����ۆ��Q����|7u&k���۵���q�mX<�7�<#�� � 6�t�f�U��Eά؃����|����1���1���=d�1H��0Q�(䜜�1���U�
�ퟲ��-z��eGdn���$\gr�*%�	��h>��,��ߪ�>��JSH����P�m�$��"�n��Ҍ�Gd�sV��9�MRǯ�-�a�G@Wܷ����:����}�&"�̗�X�$g:���l�@ֺE����4���i���c$�d������ܿ$���>��	�^���A�`A��эPL��H~���ٸ˻0<m������ot�p= �+�)`��'ӵ�Vz��;-])YZ�p���7gi:��:������-�=��&qcFZM����{�i��|ĳ*���r���qf95�s��*�2��I��f�]��@�c3��+*��Z�l��K��YY����^h�Sg�&y�g��`\&�.�X����\Z���I�tjI�5�]�Y�� 1+,�u����6�)_��x+z�� ?�x����o9�b�P����U���&����2�>��|�Ze�6"N�����3�ɧ.����6?j�S�WY��0�á��姫y%bT�P�=,���F=N/ʄPsL0�s��]vo_��w<ٗ����UA�ޣO�{�vy��\-NT��0�B?�2����)�+��z�:=�Z�k8��W�c�9�&��f�@5V�P{K$�7*N&R���z��d
���P)=yV�aҶaZ�&T:x�ࣉ��]c�d�|#Ť^K��Z��Ҿ���F~�E@l�>G�x�^� �#M6����1nPRYF"]A^&	�N,K�=_2Aw�T�`��,�_�ڰ!%�U }J�|��U�ەqX�{}�K��/tJ�o����R@t��p��x���5���ﯤ;���*@Ϊ����D+Na��~�N��ҧ �G��Kµa��s4!i���[�7��5���噞��S?�|�d�Y2�g2��mz}\tC����t�8�c�0�h
�f�#bq�@P�~2#$6�o�3J�1ނ�5�/��C���`\N�Vt̸8s��9��
�{M�־}b��b�(�����( �w�r'�_�D����hZ��w})�Q��ET�T�$�?�8��ȹ������T;}<����m+	E���1~Y��T�F����5��b��@_u���f�mG����%����������1B��vZ�?d� Ș���|���t. �I����;��É�^l3O(�Z�ݜ0�ms�!�̊n2���D�z=�*�gC�i���/�2�#`>�γp���� eK��?�
8�j�^�=���7}W·�@���R}�@FKxې���s*uW���{�wbb5�C'$��)嘑��g��sz��ֿO�zR.M�h<��<��YQh�gN�!!�m?���}�[�<�0gv&1F!��%�q�ulUrM�����I!
t��p-���p��g@���A�uӡ��k�T8�?ƭ�Sc�4an��N	����=�C�E"����}��J�SHk����	�(�����&H�1D���|Ǳ����P4p�2�O�^���L�2�؛��-�{h�(��}0�)vQ?�aF�K���Sqc�a�+�9/e&���L�ҳ���G��zJ5��n�x�~�v�����b�,H�4�m2����d���ҿvs�-t{�.��j�<F�F6)k���F���$��!߉a�VǺ��Zs�B��"��^ᮥ�?��j�#�}�t�����?XSI{z,�'�ԑ_��8Kޠ��hy"�d���+��	@1K����F`��B��x��f�h��z�-ŝ�e=��yN�$�Ҁ�/Gգ���$d�vw��5��1���9Cxw\������Ϛ^�a��yR���dr���G�ɸs�N@��<���� z�W��'�zg9�9�7{�S�c��	9
����R���f%�#��wRԍ�W͐���ا}U}`�"{�S �Q3��M�I��mf�����Ȳ~4��5��jf2��V����0�!>a0y}�C���Cqę�b��Mߊ�i~�vo���<��Q�
MW�绘J�j�L��lQ_lob>�ֆu��J���)-��T�A���=�Uݷ�<�=}��Q���f&%���a	��2S��M��t< ������ V�Wz�Z9�4p�N�nw���b{ewLl�+���~�xLi��J�~}m�NR�M��Ѷ�q5�<>��h�B�6��Z��X�o;��|�\��E��N�����+oV	�x@.���~`iP���������>hB�G���@�����Bt�u���L^�1[��*��������`iˬ�9���{�*���G�,󉦮� �q��b?{U
Nڀ8S?��s�\j���+S�.����H�םז2���f�G�{��-?n���2O�qUcuK���W����D:����t�j���\*+�P��6.~��[0Z8m]J���O�9S�}�yYXyZ�|I�/kT!��T��+x�㓗a߭��ʤ�)��G/rp~��X�pUa4e O���+\e�y~����}��"7O`�A���`���b����NKq8���Wƌ����,���� ����Ux^< Hn(��6D�u���6W'�p� �{�?!�Y�x-��/2WM�f�m#�ظf4]�gq�.>(1�g01��?C��.�<ҳ|p�_'�מ����e�E�$E�Ee��,9a�����a� `�@g��~�m[,V�2� `ro`�)p�8��8�Cy�	� �*v�nh|&��]��kc�w��EToNx���L���h5�t]�ۂ�5Ʃ��ᆖ�d���qL�?6���x�3��촔Ak�$�������8���WX�Pp%:���b�8���]�M i��f����'gI�տ1�	z;�s�^�G�5>4��Ƽl��Ń���6����vb鴓��Mqo�ߊN�<t���}z%��s~��P��@&�[���-	^�$N�펯$rχP�s�d��Ҵ=n���ܵ}��y�����%�8�]�\A��~
Kk�=_���E����3��6q'��p���l�Nc��.��[
Xl1f>��ҴR�9� ~�k��N��� �Û(]����Pjz��w��B~�I�-��]o��.���M��=�7�2W�!7#��ϔ��ua?�8�U�������sg/���N�I��GQ���g����C�! Ԩ����z�9�����9�R�����;\Xҭ�l��9�N����ϸ^*v|�v/�VuC��X[�4�S4p+��J!a��ߎ���+Z���C��: ]_?zYW��ȱS�(�ͽ�
7�<���y�
���c�i����؁�Y�d��SǼ<���)�P�h;b� Ή����Zڇ����٫�48H��˿�1�詞m����v1*O݇w�,��>�4��s�=���AI��+����0�0��ⷽ3�屚�Sɑ21dV��[�����
G��5�l|C I
5u���M�R&=��o�sQ�R��mD��K��Qxl���Y(_au�8\9�~�7����A�Ĵ����ő�-�+\iQF_�nD�=��b�C��S�>mLoY����|J	ON�\�0^�����*˛|��	Ym|��E�S����-�~���M����h�5�� �Pt�?�l����W��P�(����QP����\�̍����o�F)'s$��P�}=��JbR��2������fo�D�n�1T��T�R��x�1�_�������]���P����([���%�k���Hw�Y����y��ľ���)�Dsbkq���U#ǧ��o�Q
�J��q��!]�=�9�g�	IE��$�6e?��g��M�p��q��w+�9�}��mf����1*w%ڻ����4��kTt�Ƣ�a8���ߏN2��gl�!яŏ6&8���nb3�6(�����:�,A�8�����x�72��O��uիC�} �{�a�XZ��(O�_��ڎ$,/r������O�8ިɨH+�s,t��Sz;3@��{<��6�=F��D m??����T��2��pZ��-q�qQ��:�W64d�7.�2�:�fkd'ujO�f�lE���ǿ�Z���"��E��'��|y��@஠��9�I�0��`:���?�q�y�M�����>=W]�C�\Ƀ �V�դ㢧oh70+�h y��nə2��P���dc8?E��������Q麡
���b/Վʾs
������$�晛�ؘ�&9���c4��R�9���|Yѝ�`O8���uB��C����?^Y�V�4_Gf;��������`c�W[&՟�d�!C���EhPn��~�ͷ���� f���!pr{X�Ԭ���E�o)����c���u\`z+H�⾜
�f�9.�C���d��߮�{F��lg����+��ب�9Wd��h#:����y��1k��	�s�<c:��M_���t�ss@�i)yD�q�"��;�Ј�$$]u5\7�dQW�Z�tQN�g��o@���a�w�DH�(�R�u6��h�O�p��~l�� ѽn�PJ�Y�8��s�1I�����s+�ʶ'`�dAEEY<%�"�5�	1�h�%s�[�n��P/$W����Y���:	�^��"����Q(t�d	���=Lϣ�
�7��q��v�čr,.�c�ϴd��5�H'`��Z���@��`8ϧ~A�s&����Ӱ���?d
3!3ь ��l��/��XE*w�]A]dt���J6]�������n��S�v���i���sɯr/�;�6�!�Q�V�@D@v�� O+��T��y�ַ��sI�n�f�_�py� 0ݳ-d`�>ѕ���٬)�i�+�����+8}E�E��zD�S����z^}��+H��=��j B-62��W2�����ђ�%{2�L����l��~+�&�<s��QH���T?I	�FI!� ��A/i��Vt|�K������mPHk�
�P�tT�g^dO�?�ف��������F��I ↂ�=S�R�ww�
�ܐt���p�I���8u�0G������F�����f�BO�3ٷb���9����wk��:����
�O9���O�X�	��t�;��/��bu��p)�Ů~��r�k<=L%	���e����
I��2I�tI�@��JQ��WH!b�@T#��rft�Ԓ���<��^����߈��d�L��h0eZ,!\	L�����M}�&��,�Bq���6���s��h�@xS��چ1X��x@*��P7��y�c��t��H��=ō�wo9��HVk1��1����E$�죣�h�]��B�� �R���A��}+���a���uR���<OS�ͶC��W�ت��A��HEYXKh�{��A��y4�lT�����EF(�l�����D���bBҬ�ʷ�<]ebP,�_=�K��������#W->����'�eܯ)G��!��5n�)5c�9?�N4$i mc(�7�<h�d���J�<��Nr��'��v�&^�q�Z��˙�r�Ѡ���6��{c��?�W��ق�:��WM(FNU���|�����'5F{�DP�)�P�g�M9&ȭ��;��U�}�;K��'�;�gD��\k��#+k�AWA�����uh��;�x�"�L�)'K�W
Y�y�x 1�k�&R=s^d*mS����[N�%�O��lu���^�Sm7���1}�����)�
5.5���y��j�&<I\r�t祠�C�Kd���I<���.�P�},��l�	�L�픫����2�j�+I�I}=�M�Z��?.����l��S�Ļ��*�{��Jz�9�^�N��d��s�whU/e ��h�
#R����q�T37���7���ҫ�:��S�F:M�
yNj��k�;XN�a9(���.'	3�;]�����=����N�-$4��A����i��M3��i��~}yBs=�<����"8'uȩ������X����lW�.	��`�&]a^\���'(���<������"�[����A��X�7��K�4���[JY7��[�לF�r���} z���#����7[h&T.��vvg5A�w������!c���W�]#�6��CJ��Cn�I�`S���:���7���f���{�+�
���-B76k�ݹ�ɺ72l~}�:�bO�tjƝ��0`[�4�̂��?Z�A�5ѣC�m@�����k���丄�h	_~HD��m,�K����v���e���\��@ 4Pc�H�0jJ6�TI�f�r�b>�"}+�-�$d1��;��e������p�V#!��6y�\&�O��|��Mǲ"BBϧ"}��.'��NcmN�١�h#��XB1�3��'�m�:�n_7�`G�Qv��2��F�*2�����́KB8p6�O՟��=�S�v�7
���@�"�-�#�<X'Kv�� �V�������I% .%bU�W�����%2#���q,�r�i
��$|b+����6u�/�^�H���bp�摽���.��عi�H�+@�� ��7����qYlW2�YO�λ��E���pt����2xG�
�O��/J�L�j�����{�V#�K<�	�@N��O����mZ��>@���+K��C�e��"^���^�/�A��M��'TM,�_f�$ߠ�p���;xI�0(���x�5��v� �iI��4r6=���@�B�)�k�lH�_�@Wi�X7�B �����!������+t���s��C��
\!�]��^
\��u�e6X���0ȱ�5P�2�w�51��]&�C�R)�Ĵw%iID	p$�d�Y<j.3\N�%�ʁ�C8W�t�794��v�}�ڗ�гp4��:���٣�|;)A:��
�OX�i*>�d]	�k��	#w0G�2�>��H�J�C�=M�ڑ��������}���#�]b��	P�-�z����\BԌ�ùk�it�!�ҼY��,�KQ0�3�d��=>e9�\����Y;���U	�2(i����7ś�~��m��7ac8��L�ǻ�҂�<�f	�;�$F��������?�C�����G;Y�5��z��%:�>�K��7{m�q��d@3�r���l"��y�W�rQ'6yu�-K���t� �5o>&l �6�˹��3p:�d��"�ҳ�N0|{��N�6���;ㇹ��s+�����;����|��uI]������?K$��w7A���=��Y�U�����-�������!X�����`r�Rs80�/�t�	uY�~a�b:Aʝ��Ϩ�x!H��9P[^�nc���J`����V�"�],�?�;���B���X��������V�Wީ���(��Tg�%��p����)|N�y��܈֓�6\z�"PiV�{[^�W�hay�@P�I<��� �cS�T���ި;��"�Jm��ح��y����_�q��ŕ*��|t��۳�{z�W���9K�Z �..�C6���`�Y��85�xm�̱]��))JdU�>�P�_2aA���W�L�uq�c~�>UE��m�*��߿��j������ʬ�̻2S~�!��f���RBcH���X�+�����5�>�F鸩�����ru篟�Uqġ<��%O��J���(�~3�[�t�h��;�Rp�b�uՁ �o��
�3�j��bL�oL�{|RS܉v��LMS?�H��	O�q[��Uuqa��8d��L�:�t>c��Ɗ��+�d��O�R�e���Yl�z����-��ޅ�F�$�ݴ �u�}����b*v�Y�oR�CL.�6/�����e P��Ftm��}	lyڼ��
Yݟ�bcT����c�;V��+g�@C��4�-���^�2����$�&��,}"�nm�����EЍi��4����v5	�M1Ak�����%`͎�ň9�0�|/b���J�(���;�ۓ�x'a�oNX��\��W%����"Ҿ�j�km�Q^��������áU�F��j�w7ե]&~l�{��K�sE�9;뇐g��댜F7? B���iynv�+-�K�p����>\~¹���Z���������+��2\���w ,Jĩ�I��wF ��q�B�����b����c�]�H]���ub(67���Rn�g|dd�O��=�N���F��~3ԡ�4�ź��l��ä��Z�b�	�F;��CjH����넧Ղ�B%CV�"�qhq��������Һ�OS�:�6��q���Q��-��l�ƃG�d��	�;-˅�G�u6�AmS���BN��JTx~"�P��P�Q��e#��O���K?��0ϰ�nh���K&�{��_���GU*�9pJP���Ͼ�{��~��K]ཟ@�)�����S��*{�����
�|KѦ1�p�)!��jA��<"˞�RV\�W��j�*&.�ae�H	����W�yxE#��挑d�C|��'����\j�[���c��#N�'%0��h����~{Z6%a��!�ŷ��4K�L�
[���D�\'�n�^�?��r I�!�MD^���:��P�g���u�v���;6�g	}�4��	�jY�e���w��cM����}�����	b7���J숓258�t(��z�>q�*ۋG����]�iO�7N�9";x�32G��XU�X���[v��@ L�ʊ!c����db���%h+TY>c�ݸ��<[�B���=�`��>o�z/�K��V�}t��9�|�R��ӛF��q���$zI��%ґ�-�0Q_K�w0T^��sB!���z,(���F��SDi�}�ؼ�������T��7R�<�a�[��Cxkfl�0�B�e#�
zKZ��,�aQ�Q;H�ܻ�Å���D��G���zǪ�}��g��z�%EN	�J�i��Hl'q���Xz�C?(��a�� ��	��8�qX�P=*�}�36H�ۦ�$g/��Ư�p.֌�����ωɧc�6������
Y���|%#Β�AH�#ۓ��hmّ�(L)`��.��o�~�j�˝ؐ�fvW^3B�+Ǆ��d�=ct�q��2C��e@����}Ք�a,�^ ��C��i�$]*��x5E�m�]A�<I���?{Yt ����{�I���MhD�L��m���b�j�kf��/Ήң �͑�UKV����B�+n��d��h�B�2ry��=�� o���4΀W�c��%e�A���L�Z#�c)9
���{Jj2�� ��-j �M'��}A_�}�v�/#����Rp'����Y�T�	%X��s�av��]XD߇9�������0��J�L7�?�ZmXC��wMz&OaI_�k�7+�_#*�AB?|�Կ�J�D[t�r�g����
��1TJN;�}�ʮ�&�a��t��W�4�A|͉�)��?;u�P���`����C�Uj�nϝֱ+G�"�~��B�+��A��4f康Q
#B�U|�_�ҜR�A6��RFr�˝�������z�9�Mu�W����nV-��I�c�9�[���R�Z��hN�lj����,h��d�)�0sc���)u�^���}�аЉ2v���Վ g`��ԍ�s����I�vj�̌��Xe�2�Ul�b�$]�������ɑ�4��cb���O��*�_���~ZQ-&��w\�Ly޸�=D��#��?z�e���,3 2�������:��(Y�*��n?��ס� � ���_=��A�����aoR�*�/`=g�"��}��!�c����p1�`#�g�q�Ҕ�C!�����9U�5T�����RP�M��F#����V�TY�,U
wGI|~D����]hx�&�jmF�FFa�硵��1�}<w�؉��O%�v$�Wo���i��:�8�(��,�FVu�#M�_͒%���+4B$tȪ��x�$�q�g�@KcZIZ��V��9߅ۢ�E��7 ���y	S�6?mD FuC'M�b�T�f���=+��)g}n�CN��^����� �a����0�w�ߧ2��9况�3�]���}��F���ܜ� ��#��}o���9�,lW� D��*N� gY�����0���K��[[ǱlN�2]l�1��:��DD�4Q����q	��yk�|����|V��0�=�����l	%W׈˕Ch]�j�����]@�s�c��Ր���&�������e�ǚ�$wh^E}~U�[n),��
*Ĥ�`�ʼ��T�� K����i4s�B�vI�=Z{��{��Q7eơ{.��lP���0&ͧח��a�)��������\��_��05�
x�9mPI�17%z/v�Xˤq�b�M$��r��9��dC \> �a�'d�?o�|WьI��{|�2T�D;+�TVB��)n;��Ƃ�-O���{�cV¾�,d��T��b	��x�!��|"���� ��]A�i[^L��ډ|�>��1&��{}D��^�Q�pb�*stU��H��g�.r��;� \��!h���	/�kd!b��n�E*�r`o�����]���	*([�b��7]@�W4�dD���(m.�gvU�C��t��IUf
)��G���;AV��Q��SY�o`�?KfEo�fa\M����:?H�7h$T�a#.:18��j���O[�L�?�㲗ݎ��K B
}���yg��^H ��#P��7���ǭ�W˻M�4�H�}e�I��ͽ7b��N�H��z��I7`����2C+��ej�_9��H�y$��2Z�)�z�n�B�>�*���7�1,�$oZ���
)p<�S4m!�S�z5�q�sK�Ѐ�/ ]/�[�p�v���f�?N"��,�Ni`��/L����R�P�}��� �E #A ��'0C:�8,�el��bz�E.XN���](�i:�}2t&9��j6z�h�W���v)�R�6���k�G�x�L�ϕ��a��������{MZ�ۆ���U*r)����8�	�4{�X?�nv��������4�x�3�[�{� p8ވ[qd�iC8�W0�d��i�y0���4N$�
<-o=���$��D`���Ԥ�v�%�ߴ��PETai�h�Ǣ�F�:_��\�R�����P|X��csT�y�(p�
�-ɰ�*1�f~ѮO�	���
3$���◢�L�P���O�H�.̴���wwu��!w4ƕ?�3�q�\-|� +��1��U|?/�q��4F�X����J*�ĉ����L~Z�w�qe���@�I�Y�"�|� !�� U��9v�g��Xŗ�c@�KC�Q�?"�Dh�Q�aj�-n
���Wi^v�a'�7�	_vħP�%sY"���g��a^nE.����� � ecq����Y�!sn`zi�G�2��*Ee��j�yI���:�̷8��Z�]Ei񠁸*A�����%���<����?�a�e�u��=^}F����?jb�x01��������kl�f��O�դD��b��"UT�yG���o+���v��%��$�6	t����g��m��3�S���~�:��Sr���g���Z<:j��8<t��Nx�ٮ�"���z��I�d��˚)�\�����?t0VG.,��
�V��)�Xaf[+��GL�����KI�%�BT���L�	Lu()a���z:��rP+���i?��)��I�k5��h]��"d��=k%�G�g�:��c�!��K_Ҕ�'(�c��.���Q��؄AF������ch��[��YʗcX���9�>n���͞G�:�e�}��)d��s`YCD� �N �~6tOb:��%�M��ؤh[�hM5n�}�����{���Op�V�Hf��Ӏ�� ��� }mV�Z���x>a<�s�G��������>�� 1�42M��a4Ӏ88�����*X�gf͉](��"�*X�S3�I����\�Lm3�2c�R�{/?��|�kL��2�J��#�KR���@���\-!
E������ ��'��c�=&l��1��P5��E@��>t�.��gR]������@���w ��bU8�p���1x�[S"���2!0n*�+�?�R��S�\��n�Fe��.�eZu_�"�����|��W�8��~������+�ޡ���l��J�^��Қ��ADEC�����VFxmGB�T=�Nk�H.ΙRX�&S�!v_����r��zN�-u؄��?�s��G-�������rd�)zԈ���z._���_��H�f61�{#5��S�W�U�L;3�[�o瞜ɔ��-��i��E���@�t��4O��{�d��O�� z�S��aQ� � VM攭�'��'8�@-���[^M��#.�d�z��co}���*�ޡ�\D��N%מ��5rhʇh��d�x����(w��r�ԅ@D�(Y׶��Q�Y�jl���ZN
��E���,3�
�����{�:@���׵�	���z����bM4�Cv�A���H��V�<�#s��Su�^�Y�.�L�Z<N)<p=�r����j�3?~��D��L�=r�L���TC"���a~:�qY�e�< T�Q	=�=]+����_�=ި�
�w%�:�]��Rrf����C2�mxw�So���f���
#:�������!
�_?2R�H�M�c�3P�!�@�u&f����93���3��<r�L�3�(�d����F#��3��p�ϡ�b�r�������dB���Mw��&�T�r㙥�J�ق����z6v�啑�r3۟�n���4�����_��A�
�]K��!����9�`>��z0���\�U�br ��n��]��g^W\>s�{����j� a�/�ƃ
J������P[Ôb�m�(�s<���(�	�Pe�y;������\_2�-��c��XV	�3���Q����)�k�P ̹����}ֱ��&6�G�2����M~⏖���]�����b���ӫ����� �5%-K�q�`Q'��(;D���Ra�
�G���d*�N��q!�!�R�OԷmz�T�=*ٶO[s�y���z
'��w�?���75[� �qJ����st����(î*��"&�0�h�<\�~J�t
��?2�|k{�QP�]�^��-�:M)Hg1�D�(���f9|����8t�f��1��M�X��2W����**aw�!�ݐ�� ��T��:ـ�eUɘ�y!vfhN+q�+�ê��G��6Y�Ĭ��pʳ)we1F�XZ�q���o7�+J8|J��y1
�F�H�p�-�
�����ط�rP�u׺X:GbN�?+��Ǵn-�R�t�r�(��J�4���1�nR�'���}�y�������D�a�&��+�β���:  �N:�m`��ԶL����P���r��R�'�s��>i��%��/���%#,��淪�o�i
�%!�1i������#>�J�LX�$X\2-�h�v��Pq���@��űC���ڒp�\`R�)�p�xo֬�������m��_��A�@Yi��al�cTq)FZ��[_N���B�Vּ��h,�o��8���{{�T��Hʚ`5$r���8-���e' �ӲI�YX���Fw\/p�����3C4�Yȉ}ͫ�R�Z�y^���ڿ��Mv�����T�GUK)C��V\���֣���@�=�[���H͚�H{���r�g�[0	?f���·g�@�(\&�#*��7�M��Oh�?[�X?2��V�Y����½=T�m(�����x����1x=�xX&���Cd�0V,����y��|"B,���K@��%$e�q1��0��:[u@7����.�I��n���(5^�"-`JR��&N���]S3�
2$���)I�璹�(C�k'���D��Y���sV��@�j=�IZ�A����n�̝�S���ڂ/v@�R��,/x��Q;�� I��UC;^I�'�^NЙ�n�4�6��K��rM������k?3�k���ﴐh�2�*a�+�X_�_g�c��E����G��'�3(���Ҫ�i���'hi*�(����U0���E6��u�G���XQ��f���p�z�_�%ȪI�v`r5����d��z{L	�����Zc�1�N� ��eL|q�.��Ĺ����r+�g���E�^]}�U3�޻���������@f*��Z;x]e����Ns�w�c_��]��6�.?��zJkc.i7^H8ޠA��k
J���3�6_������`��M6�4�Җ�����?�/.���	o��8>�D4Ɍ)\+OL�����3@eg	��[q�$a���!8Ѥ�,mknL �+Uk[	�M��`����/�#6�_�gDN���B���EŊ��rP��m�s}$��M%ق�䢃{\�:td^��Wc=�m��#����aQ�T}���z�@��U�������-.���B?�����i&���M��1�����[���@ݜ�ὑ���ߒ;�$A`��i����8�6��q��[��S����,8���N����G5�6r�(�n���$�H/�$!�����&�� ��%��F{���&��"<��c�$-[ �\�!���'A�6���G�U,�C>��HABoH�ǅl����X�PS��Յ�{���s.<����i�֖o!�E�m��rњK��l�[�9�Ku "v�!�w��k)���m@9t�Ua��lo1�5�X���9��i_W�Y�;��x}�x}A��>�Q^���7eH�lK�IS���������V�B��q}��n�ԧj�m1�0ܤ�Q6�c3��?�}�=1x��B�;4}����^̗$}F���ad�x�,*���Q|#�Y*m�j���ԙv��$�9�E~*���I�1����>����'�;3���S�w{�sA�o�߻�C?��~��k���j���8WŤR�0��rH���fJ�u	{�ǻ��wpsʅ��yO��P��n�П������r���M�⠆��LGK8�P�5� ���WV D�|����s��9�@�}�%�M���� X��]%���U8t�k��y#e��,ki��h-*Wj	\�l9g:�XY��/��� �B��,���ǋm�N�пpǌ��҆4H��s{ �n������}a��V�+(��C Y��i�Z�� �p��ؿ��w��,��.򷈞0S��wg�󟥀�lp)����z��Mt�hb��`���X�%u�%j��pm�A��IGǱ��|��;��*�!VѐI��{���5B���bRJ��vxp�k7a�V���`�*5�Rw�F#�MN�²Q�r�ib�G��
�'X�䂱N��݇�6��L!�8���r������T�t�mU��" �����S�^�!�-�뷜�Ҷu����<�[Z��u�f���A���2r��;X:�?����hC*��tj�|hk�z��$�Ix�1��$ǔ�T�^^a"�b=��l�eK�Pr�k�����R��L�f�EP2 ��~a����{�Po�L%�U���-��qu����^ƶն������v[U��3Z�����K�r 98�`Ф����Q��[�A�^6F!���Ҷ�@������T�ش]t���Յ&�)V�@�(@�+H&�ei��O i��9�$O�=��a�.�G�p�9��Ș%3Z���3�&GF�eW�f�R�gR#�{84��3шVKH�H.݃iҧKI��Ժ��+���u)H���~�4�����&��{�:z��U�!.� �j7Ј�D�t�k��xhT�0g�����M��GƎcߴ�X9���4S�q�ٖz��e4�Uߦ�eu��Χ���P5���sb�r9$����(�ca�Ύ����"���Լ���B@}.h�^�%;��P�1��7�D�jI�Cf�:����!fLϮ���8 �p�Z�fa��H�� '?�.&�X=��B�� ��s��Q���ĀU;:��<��f��6���Q�nn��H0Pn��������	e�cSu�C���&r�r3��m��F�$C|7>�4�ŵ���Vħ�NO�}6�����:M�D۸��/ ȑ�娖/� {꺘�ۏɵW�mwi��;��X�A��dM�Ea![Ubd8G�-LP�-\�o�k���B�t�Zi�~"��A�����6�@V�r�΍/�"���Q����;��ވ4��w�ck�g��Ē��;�J���kʤ{����)�񢥀%]"4�*�%��`�9B/߬ĂH��s�����j�W<,Y�\�&��{Z6��j=7_��W�7��I�d�v4Bt�iJ�-��=�M�S����bM\���-�#�w�`)�2ج\F��z�y���/�FmG�r��w�s�P��<oproʘ�я��d�C��������dJE�ͦ�8=;''O7eN�ɦpj*{���fb���_�j�x�����zG�8�e��c-���(��J�#��"5*vq$ p�o�Ho:���TB�,d,�h$᥊��X��@�aG��rZ�T��#����S�K��+lN\�ԁ�A��Df܅I�L��š�1s=�|�I�@������NJ���\t��̬�^�2�y�,{kNw�ѣ�9soV�I}��a��H��.�&{o��������an��5(�x��qҁ�Lܣ�rs��,�������3�fߒ��%�䔴)�é�6�H� C�S9����-�\W?�h��D�,��7�1���Q�y��a�fs���U��l�_7���x��2�����:skDZ��y�!_��J1rM�6�d'Q��W��isR��}���K�P&���}YB�>���M�J��k�<�B��j�ݺ8gWf��d�'�>�1�/+�!/�@,O� �j95A���S���-!_�]G!��"����v~��,o���&|�ۑ�4��c��p�ky�\����P@rnG]�.��m�0���A��13+D.����FȚ&os�����k[��b!]�$� ��s���1r����ma�Z�^+X�҄��sL�g=���9o��@IO�"����տ2���L��hAˍɖ���x���Rc�~��=xej�j�=7�,_xK�"��W�cZiQߨ ��І�@��� mK��ȍV�Ja8Ma�T������.xp�JT��^�G.yDq�����fóq�2�eec��+��+_3./�]+ �ӟ@/E��x7���ˑ΂$�0<�60���s���l�53���E�`5��h����_+��U��B/;�}'���6�$�G1�β�h�͐eS�B�>	�+�7d ��'*i�=m��d�y��O�⣊�;��4c�^�Q�n��u���΄��8x4ҏ4���~�d��+���]U�)� `"��[Xy�h�%��!��V	��uwE}s�Ȓ���a�I����.�~D8�����q�t��,)0fP�X��/��{�gA�s>,`|B_�H����T,�ws��Q�4���T_��!$AI���3���TlX�@�,W6ϴ��ڒ�+.@����d]�F@���eni}�UF��V�Z8�� +M=����r�I��QT�D\ /͓͐Q�*��yz)4f��	��-i.�2M��فM�ק��+Ǎ[�>
yv����)��y_*��g����D&�l�D���+=D��<�#,g��3�ei��O6g8�x,	�=�	�
 yMT��(U��U�7��ٙ��T�9��%i/e�2�L^�jc��%����0��#�0"��P�Rc�-ʵ�LV���Ub�t��zekƉ,�Fn����Qŀ��,��1AJ���)��8�h̎`�a_a�R��i2E�!Wg*ߊ~��QP0�T�xJ����+�]�%2�C����:�DȚ�G�n���DPlB��d��'3���$+�c�}3.���������U1�K�R0B&|�]�㖅-���^���6����NpG��ns,k��vb�m6|�{�R�"�橰mB�w}��W��(��%���:���"��Ir��O�	^��B��ad,���݋/:�t�
�}eh�A�ç�D�R"ߏ���<�S�LR�P�g�i�p����qj1{����C~�G���w+�2���ٚ:=Nn.�Ԭ�o�(�HB��(ꈩP_m�|�֩s6��3 �{���r����ώ�q�#�VJ��	����>T����6(y���}���#�R����n�v|îwt��~�W����R�E�]S����@h���1�g�IH/͓��4'P��s�)�� #w��g5�F��<\%�N�����x|jeCՠ0�rC	b�mj��*����_�3U�?
�8X0�NGN�TͦVP@��vf��~�$B%���CX��"a�pT3�e�
�� �3�G�3٣�Q��H��C���0ޞ4�oq?��8ey��oDVkT#1f6�+D�g�VT�o-a���YDo6X�D��bqvf��S�1�U�X�˰����	E�2��w8��}w"���Oy��]+���Ѯ9�c���(.���C�ұkQ���=&� rS��h�~M��i|���xH�yt��3�����(��D�bR�q���|�gM�%	��*W�*��@�/0t�"mSj4ЫU\Vq}���Q0X&�ˇ7��c�$%���M	6[s����xm^_]Nv��L��6��1T�ֵS&�����I�	R��B����~.k��YP����Mo��Ԙ�済	i}"x��5H�,�}>/��X`)ryz���6.v��N&P��C�P����[K�ClcQ݈��$�K�3�9%��tX�/Yz��'Ը�7V�NGs�-|g��IR~xOo�Zu�Li�Џ����ҙ۠-���}���Z �5� ��j|4Q|�O?��+����D�&����&�e�*e��K9��Q�+L�Ҙ�?�Ra`�u�+E�3���ĳ��L���nm�)��$���.�ݽ�Y ���s� ��?&�WC��D8�%�=Qp�2:�RЊXy���#\S�S�&��$IE�Lrk���b�j:{QUt��z*���#��7�6�]'	���/9뒈"f��c}y�}T�`��>K8E�I��-���ƥ7��k��a�$80@�f�����nZS�iEk�B�B=n+U��DC������b����q��$t�D�	�SZ�7[*�ᯫ<�!���z�L8���}�j:����������0կ���N����'��*���������&i�@����@�5������"�j]���r.4��Gfk�r
��ϛ¼�v�G:�����3�M�Ghd�u#3ʾ���/�v�tWgV�TF��
�YBWN�r��nmr�vĊ[%��D&\��-�Q�G=�:mA� Zky�O�mD�d0��w2ٰ&���l�&�rE��^�5��\�� >��P�=7�&�V��Ѡ���mX�4����U�ҥ�0�#�JU��8�꡶�� �zD�he�ݫ�NR�r}Y�v������b��ED�f�j�q����A} D�T��.yb�#�b
+��8���ug(�՛��)đ˹]�����%�*sz+m>�d�<�ժr��`�`6$��53��+�xޓ�1ԥ&����ux��.�N2���O1��^"��_�0�vG�Z�0㵇��զ"����]�ANb�t��܎.��5ow܂ZD
�D��d�t�˾ۅ�Kz0ı:�uO��憞���ס7��HA~�R��iM�$�^���3wp�9�_|�߃�^�=�&e�qj����/�f/���	ګ�rŵr���Ƙ���M�4F�����&��\\���,&�^�w{�����_��4�*Zdzْ���/���Bxp�wf�N���N�~��ػQ���sUp�/���Z9l�kom�26���G>(d�Gh�B!�p�%��h&-�k���܀�MW�r ���a�m��h)���J���햃7<]����I��]b1�8L��D^���B���x�g䱽2�$���9��!�2��u0�G ٲ� MY�wLhBP'���H����|�i
�f�߯����H�6�p.(X��Y��(!�Q��_�Cg�Rt�J��ԓQ����'DS����6
aC�UY�6�@�����~A�x�U}N^���Xn���҇��zp�R�&"��'�gS�k�Č���ڜ�u%8�
љ��ַ␋��X2H�[�R��]�f0�y������W�:�Z�LWj�@֘e�{��	���,����s`�S$���V�����yE�A���Z.�3���2�T�Źkk�,�xmm&A�[�֗���9�1Z?�iD��ڋ��G�:��"�م:��qH������L� �P�㿚�U�>!�t��9�@0����M��e1XrG$
8ޤ&r�_=�k�+BZ�`��3ִ�O��+��Z��-c_�Gϕ~GO�� 3]i�ybϪ�hqב>�
@) �K����vu'��nGK�>����l�.�
��[I�0`;
�D��$s���?�fn	��~�Ns��*-�=�]~�V B�-��
Mh>�{�V]R��	
�+�*w Bp���=�)���M��_|�R�ʦϨ��1�kt�� KY*�D��`^�����t}�'���+�-p(��)0|[�Zfy;Uk�a��Z�}r�\�djl�O�>�X������XwK����<t�x�u�MAsԋ(ǣ�O|ϗ�S9���C��y((9��RN��S�;^�:	v��W��di��)�
S�*�����緸~Kc	��xvGpa�g��R �i�-���w�
���m�ei��h;� ��� `iDS�&�G�Mh5�)����|@奁�.�ٽO?@�a	�@rS(,��{�*%چ�n";e���D�[JЬ���QCUh�$>���L�����VܥN` �.�F%__̅�%���J�Cv��a���֟��ܼG�3U�q�0����"���{~��t;@{i�ݵh� �4h"����C�׶P��p����j���c������H�_����9l�����ǅ�V������a?�8{���}���/�K�G����$X�����L���3I��`��(��Tpe�B��h�E x��@@�R�{��Q�g)�:3ww�p�䄠mD67�Ds$}D��z�k�@�P�,=�cT~ؿ�B���b�w3LȤm��f�<l��j�h�40s�r[1yv*U���<pN��O��e28�%���u���z����m�Df�[�Bb&2I����ّ9��>�LL��(*1ϰ�w�G?՜��1�4�����׊�`TS[9!U�-��#a���]�[��2�B]��� 噠�T��{�ʴ��w_A�~Mh��e5�˻�R�b_;�����
�CG����}�4����>��l�w�(��ڤm5{Vm��
t��ť����Œ+@#,cd��b�;I��C��?�P�q#��o�7�q�{��=�7�a^{f�D�O8�O��%�/�sc���̕MȜ�0@>�;���1,���H��j~q��~
6�c͔���,1ۇ�!ر��9�%�v��YLd���j*>� 7���6�8J��1������8�z�k5w�z��q�M��Ux���vp,[���^�x0�14� D�%Cn�̎��j��)l�&/�:������ {(Z2��xC�Ie))�߈��ۍakv�!��Q��.��^�^c�:^�_+�k
�wq�)n�@�`D*�K)����",W�?����Fk���"�8���:/:�"���#	�y�w��G_�K��q9� #;�*�6�5)[����8#uR(�ڗ��__;�y�I��^G����f���TZX�&��R�onƙ�W���j�P��!x��
�1�j7�yc����C^��Ϯ�����ieβ����ې���ω���JF`�N�k���m�6�^Ǜ��t��V���<k���'�z0��d<IS,Հ^ׅ����&����̹n2F|��!u���U��q�������t�k���1�q��?Q\e��"e=&Q�r�����c��}�M��D�Xc��*[s���o�>>�����[��6���LH�?��}���Q,:�sN��@��)b�� ��Ovݒ?�Z&*,�bJ�D��6�Zf��ߙD{���t�(�a�-a֗7�������[���t�d".�N��(��.E.�ce�kb�����1e�4'C�S��qE����q���
p�r�8Z3l�UC<�ȣf���@M�|�����./�vMu0�~�8\���1�����z�B0\+�������|����[�(úC�F��- �ɀ�I`o��]Ć��|�4\��ܜ��1bGPG�
� ;'
�f�}<�����ʏH�E���7��k��F �'^��:��u� �(�R�Y�y��a>c����7!Y�^��e��z����ï���2燯?��W!�tO0N�f��)K��W[�-�㧌R�� �
�����'���y	zKQh\��`T�`͕*y�����k0��֗j�F0��Ǐ��	��N�+��V^�~�dt�6G���1��nS6�z*X��~`��1ü��m�:X��6�YJ���v��eCB�%�.���3����P#�i��A4���`"�DTT�p�  e"�r��VP����oӰ�n�J1M���v��U���aa��ߖ^�4��{��)�ȀeXS�?J���a|x���7x�t�$���d�v��𧖤s��Ԛ�s.~�@�"hN���W����L�5��i�
"~($t��;�=�k��L�	*�4�pQ�ұ%��2R�ˏ3�X+���BM)��:�ȥ�oB'7���+��) �n�,�W�d�����Q0v�ʈ�����iL�Y�D
��i�����l�K	�9 t���+�܀�7���?3����6}���u�E�:��������@|�G��B� ����Yfq�����y����CȲ�01���Y��&�/a/μK{�F���?,��߫���'�X�&/�\�p�eNp�~���T&�?)t[B�gf
�)�.I�>t�;����\�gI�C;�@$\�d�)���n�a_*����x�9n��iZ�b�p��u���!��tɥ�����9uk���}�>�s�ڙ2{�m�Pf	���1r�B1�3��2E��Uo3�gu뮑�dSm��Dge�a�%'�ISxj�{<���j�G�=��nPli��%��j�|�N�DϯL���;�t����q� v�-�����2��B*ˑ�����a�~�O_�HВ�d� �4pIQ�t�������~��ƚ�b5g��I��\efT����M�~�zj��[V�=��=�t�����	�Pj��_���ɾ6O�[Lp���J�s�X7����e*�0w���'�%�]1K�^�ma��`��#�O����[��Z�{�� �怖�ǁ1$�5���Y�^�-+r�Q��R`7���d4�)5��'�)����^\��Ʋ�T9_T���d.�L/�4�"X����K���Xm��0ʖo��J��^��o���H=�+:+�k����O�u�a���j	���.ژ׉$۞DH &z�>�6��b��FX{�@�_�N�OW�f���0Ik�4�jlqjV���f��r�\��!��;����=P@��˒P�o�,�Y��L��=5�݃(�1��i�k_$�4i���U�[p�v�!�HNSI�$���d���׳^:u��3����4�W���ɖiB�r�?��*[�-�a�\��,�7N���gE��,MU}L��Ӿ
�>+�9B4 �f}"l.���J�F
�FW��^)b֛	v`�!�����{���W&�Pǐ@ZD�CI�q��`L �Y�H~r�����K��wF`MI��9k�QJ�^Cr�]:B��Jr�lq�zV��oq:�B�S�YR��_�RvU����c�~���8�G���Yaa���[��5��Y����㪦�7�)��3@*�[yxr�6� 9��j��@{�4�����z ��J. ��ˇ&MD݈ /�YǣWݯ�OH��ĕL��@�E��x�RW)'���7�Y_{�2Ғ��)˦麤'v�@��֒QC���rG �y"�/�x�������z����u�$��0�I��	[[Ʒ�A�lR��;����J2#h9ٖ��Jو?�{Y"+kt #-NcW��!A�h���	�rM����gD��ˬ���y���,�̨�k\p��t�ݞ]�y^�^Ez�`!h�E�~��fǆ���q��%���&Q�N�|�Y˰�L�E��OV��[�$AD�����32�fԐ:
�}�g�dB�jM����u{~[#!�I|��wk#�M�%��C�V�8��2��Ez$���0:c�m��@�ػ�� g������%jWO��J�@ � ���҃�0N�h����J&_&
(�@̗h�	��^�u6U��-��&�uE���H���P�����A4��yh�@p7���������FV���*��CL`����=�(y|�
�uc�O�*r[V�=�IQs-֊��C�\���n �z����,]�G�AO5	�:���q?޿�O*��r�l蛚��y:��ö�b�]�4���3�4�8"F��{{�o��Q�C�0Q�����6x�_�j|����-���Pӑ݈�Wo��(�K��_*��#D5,{Sg���~WR*�h��{�Vt��� �����	�U�q�$��4U,7[�@��A{ML���	RNE��`�/�OkxP�(�]�|��|V+䐤�hA��(��0I��8Q�F�d1�IIIjt��T-�葾�/H]���g���$m���K(�֖�ŕ����x�A�V�0a��m�*P�'NwSN�N02ў��� �rSaG��$0�77��x��� L�.��=��O �����$����ؿçj�
K;IJ�y,ti$�3�b����xo��Il$�ClHH^��Y�QMI3/�(BZ̻��5+R�]sMr5���SzBh���@�����v�a a�ϖ'AQ�,f����無*up�Ԁv8\� ��v��>��uz����)��� ���I�"�_d�V؎`_���4�RYX9V��f�п�	%�����3J�I���l�qh�&�$PN��Ʀ�������&��8�Hپ��Ҽ�E�>���U�t�Ū������ɜ�Ϭ��vA�Y��~�v�'������(�������:�DvD��i��]���N�/R7���o�j�#���d�*q�"s�����
��[B,�t��01�ÆN�m�!�#rJ �K>�Q�v-�4�Sc �i=���3�)�C�CBŏ|@�Ah���b�����M��N�+%ʑ�����r9��q�hr0�M�w�:��4�R�MTPH���гe�^a������$�R !��i�-��zꍌHFN�����cb��m����'��Yh�\�Q)�6��o����cX�,�U�����i�'�g�1G��#���2�X5�V
�L��R��^�����OR��1㿀�B���{��ĺ�y:񧢹g�ث��%�<Q�8����T��̕t�3	V�^ @�2Ȁ0Ht5��vt���(Y:���&n�z���Vg0tK�� ��P��'~�n�>����^V���P`2^	�hp�=E^�5`��K喀�:)�|"��c�wfԔ���,w��(�N�a��\��ξ^��]v���Ywr2���E��[�}zFcɠ�\�
��sT�}��ӯF<�5����w��i�����w1y�50��>��O��`������R���7j��dT�;�Z9R��vPĈ�X�SK����k����mB��p�u*-@���[�_�����p�R[Ym?R��']��
>/�Ben,�r�I�/���9��O�(��E.α0�Js�͈������ 1X��tM=���y^���'RS.�*��IڃǩSʋ���61�'��|�*�c�+��:����H����>U�F��")^�[6_y�+�������
˝�j�i`ݟ�_	���{�fN}����^ǡ�<���/���M��	�w��]���6Ʉ��M�.(,����]F��1����n�}b^XX�|B�Qh��æ�tQ(W�,G:?��8A#��en��a��@$�v�3�I�:�H��G+[q$M�yל����!�K�:P5$�D�
�hOt2����Dv�u��G]�:d�,O�~LX��I�%��5�{��BTX�,�N�)��΂�1U��;o��{}Z����S[N6Ԭ��a2v���א��m�.�Q����PP���z3'\��"��4�Ԩ�_ �qgrXdGvH��BL|IJ��岫t�!h�;dYBvP���w��ƿ�(*�K�7��tOn�/�Ѕ̌oQLr<^�oC+q���%U����"���޳�գ/KU�xN�h��$��,��*��|���k�|?��!ϲ��F"*���ےZ'-f0��?	�ɪ�_pZ�b��l���N�hr���Kg��3Q|?9k��y�+{P��ǲ���|�y���m����-�6��5���� ��E�k���_�3�[��jS�:<e7�	^sx�S"}7��}-W,a�V#�a6�|�?Ɋ�[��$+�Lu �8R������~��8b��y�WkC5���3�fv[�����uJ."�0{�*I34@]�yz������s�gk�ɂ|����b[�."5��mN������>Q'Mu�Ma����ES������h�l�㕍��=	(�n��X#�""��������J �|H9�g�v�k�f����H#I6{�:�b>`�,�����X�`z�:u��eP �L�;u�������lU��-}E�{^���� ���r椭yl��{��)Dp���*�yM~�^�s��ċ��C���d����Ժv�Y�Nm��Vq�{Ƈ�E�g�,#�D��U��������B���mw��H�,}:��,�C�9�:��Y���o�:(H�zAoM���V�z4�}_>�����:p���.��ນ����X���j`�d�{��˒���d�b�Ť�l��gn�/���xI��2��Έ���#�B6E�6i�y�ZKU$�-�@1j�B���C�����;�&�u�����s#��Em�lOb��@�̔�̬�h#��ڻ<h�Tn��S1{1!cQ8�.Ӊ0|3�Z���P���͢��D��e�A
�7Z.����9������3�i�\k|ֹp�����J�'��!K��`�D.W%��7��1��Ц=����l`���Q��'�E�$a;q9~i�n��`@Q���X(nRv��,'V����jjYAM��L"����J2���v3��VP�*��/B�MS�y�����!���;�H���|d>���R�Jg�B"�$Y��yN�w�M���U�^�b̀X�U��H>k�:�F�s6���>[�UQS�U�8�n3���`��q�f������������
'���٫�
�j?�ǻVQ�G	�r�:�DG�`���Ki�Y����z�|����9Gh��x��.{c�l�kŝŴ�E���������uC�Sww&���m�9��7j�;��T��<���G�[�6T��=��22l� �5�p�e�'b � K;BX���(���Э��&��ۥ���/��� ؛8}���^'c$����\5���)�'A[�<P�ܸI_?�����h2&�** �i0�$B�.0�e�R����([��j�-Z�{��i&�N���SČ| ^Њ����?�+�8�g=��
�mƏ^aϪ�ɞ�12��[Je!ϕ˧�Gz��}��u5S��n��;��RO���_�j��r��)�vO���c��6(A���"j��c��o��J[l��i-�)�(������,�ބ��)�Q����";[����>)�j�����9�Ƞ�&P���wV��̴��	�?MJM26�Rad�}BH_�����,]Rq�_�u���B��]9V���GA���mxV^4��ww/0c�M��!ͅ�gұbMɑ��ޡ�0�s����zZ��+����@���V���O돐�`�d"��)m������b� 7Xb��	�`��q���U�ʞ,�/��u� M[��4�_�dm�O���+�����α�ۉ��%��b0��=Y�{�D�� �8Ҽ4'�� [N�S��.M!�6Ԩh���4氂����	|ǚI�A6=1L-}�+��KXx5�<΍��>ZUvY��_yg�@�&�2�rLiz���WH��]�haV/�;���>vW������	,a�����\������T������h7��V��
�xE�'��U���3
W!�5� �G�;Jh�b�y;x�+'l���A�,}Z�F��H��m� ����ȗz�wt1�jKKeW�<"�A��{�e���l��Dш0q��BZ�wR����Ye��W0:�u[F a/u�Vॣ}Z	��$+��Խ�u���s����3]��ڈ����F�W�Z���Z�����	Ry,QִvhzX�,V�g[M�΅W��-y2`�MNn/
;�*d������GK�����RCZ�]�_)W�����3,�½��Y�-���3���V].�kYY^����Q�$]��i���4�E��A��>�G ��GDe��ް/Yv�a_Q*`&BT{Q&P���M�z�/<�s������[)qZU�~�x�����jZ�7�ʣ%T�8	����5O�,ye ď�����2U�u+�X��2�<�#�h}�=��<���/�+'
���u���8;�����oz�f׃N���3�d��~��K�w�y�	8���s��Έ���?hqU;�ju ��*p�0^���(a����%���:Ę1.ϰ�����Ó�����u��z�ݺ۵�o�\��j��Xd]4�z!��ǥd��^Q�U�,::���<Y��,�l�H���� |XCH������|~�c��x�[��ԏ��sV�ʧ�_�r���F'��qt�4&�\7�K��\�6��F��s��i�T�ɭ���-e�=�t�,�	�eZP�G�X[,6���͚|W�����<É&�
��� LM�87��9;m$0�O�e��A�(��j|W��!Ȇ���D~IaB��^�	 ��i��4�)�?2��)�^&;��H�s0l9�ϜŚɎR7�`_G�@����o���=:�wn�ۜ,��Gy{�v���X�o=�iv�O��Ш(�TZ�L7�l�7�.�3-�@�j�u�jx鑓~N��,���ʀ����b����DWN��̴S �F�e�p�,�1��9[_��y���UT�`7Zf)w���p��`/z�^���;�yc`�*G�f�x�ғhZe����)�����^I|G�{(���>�}��t*��\�:;�Ӟ�s3��̕ׁ��%�<�0"���#�I�
�V\z��Y��;�?���hϣ�[C.W��z@�r ���Z]�H Z���H��$.3��V��_��56{��w�iFY�E8�I�`X D�Wiձ�G_I��y}kS�P*�q[ߙ_�����D��RaN�ܙ���;ۛ���J�������K��_i�f��%�	eg~c@dH�;{-l��r^L0ounb��l�ǫvF��ݤ)��"X�I�T9��jLɍ*���7������|~�q:��-�Z��k��X�9��%K�s�`-�{�da�g�՝���}ֲ�#�$xY���Gz�W
H���1��b������C�C6-Lg=����p7l��NӞ�P�E����h�/�Y�2��+�T9��֩[�F�0��_�&P����9Z �0n&�{� gG0ӽAD���ЧL��z�H���gdn��V��[�[�r~��u
1D���O�sƔ���yː��b^�ߤ���_�  �E�R��kz]�U���5�j�9�����,�;�1�1���U��RbM�M��?��H7��
�h�K׺��r<�C�^N��>�[�w�<u9yI׹eU��H+�ǣ6��mP�v�~�g�X]̚�����O6j���:'�]4��s��_�#r�6E��ڄ��#����焲�DW~h%��0�tPD�1��.3#xY-��3��X%�Fw�`8��mss8tp(��RR
M�����iLu��!�8Q?R�M�z��v��A6�dE"e��.�TU�1�^;��g�����='�H�=3�&~�|��F�i��.�L�AQ�^ l�Ö�W<���Oh.T8A���E�X��O1�Zd��%5֧�\���&�� ˍjf�sJ�I3�g� �ۇd���C���6�D��b���{��a��"ND�GMN���4@�v�č�{������2ɻ-hL�7�<E5�M��a�f�ED���M��>C�����Ã�RB�����~J!j���>�A��&zxA�-]e
�=��j&�8��y��6w��w1��?���2�0-��л�g��{�`��M��w�4�}��,��@����B4|�������'�L\6�V��x��"y��\#M�v�Ve%�ڗe�Y�Ѕ� Hٮi"���(��q�>�ٲ�Tv���[Wk����W?�ACZ���x֧���D�j�!ત��~���h�="�#I.���x�e��%�93��բ�s���n��p�#��a~�`��p��쁘�tcɩ������_+t�
��d�pDU��O�/�.�y	z��E�)'Yh�0���9����ͪ\I<��r"��l�:�@������-���2b\�j���3~��j�~�&���_/�����[��K+fќp��� �S@g��1"�"B�5D�nL�8�Z���;��n�4�1N\q,#���G��_�Q�]�������"h���l�	�<5p�*�h�o�Eǳv������f��"��(�7��|�âgp��K_3=���K�zʡ�6%n�pk3X������-������O[z�y1 f�H�p�d����)�p���l��v
c'6\ow�ّm��?���� X9�\Lx�B�*�
�^��:U~�����w5S�@�^iћh��`ͨ���!��͜�
e?��K����4��N.�͐M�<�\��]�\ę�m�s��V"�M\a��T�m̴��묾���^�/�#��WL��4��Ē��l��U�eqdE���~^���H+��΅�gp�^:-G��VV�#��q(�́���D�9�h}�3r�S4:�L�ʝ��y�⶛o*��ͦ�Z������l�i�e�1Q�8���,3��<u�M��י���z��/{���q�������aLKGmΧvP**�X�
e��#�*�YkP��P�b��[g&e�-���$\d�Mo�>(aQ�&�Ӑ͜�C��^\�*F��x�� ���϶I��t�e��Z��tL�+��%B|�_��H_7�->G������cÅ���Dk0)c��ьI�xq�/@�ֈ�y ��<{���=iP�up;2<�9�� N0�m�l҅˅ �`�	]��_�4A��,dn0X8�{��\$H�[�XG�kF���=�i�X�3��7�c�jJy��3�,��Ƥ�q���<8�/ͫx4��:�[��V��l��~�?�ix�>����`t�b�a�f�6�.��A��@�]�K�e4_4�@��^R��{��%��_NDR˕mm�p�o'j\L1E(�'I�1�'���O15Bm���Vkm$�����d8�w>�u������(@5\KD`�T��/�Q�����dW�0
ў���6T��5߆4��:l���mi��LWE�-�GE��j�n�~��O�(3�1� <OCa�}XnF��=J
�h�ȿ��	����vz�����B��H�i�����G��,�sq�h��A��ν\`��t;z�u�]�����O�j���3Ҁ�x��·]����;�m�$S3�ɹ(m=�(l]�x5V1����&6�JH�C�._�^L�/j���S?��p�ao]���Ls%Rv*9�B�;0�]�J��7ݥ�����Bv����%��D'\nۼz�r��R���!�Mګ�W���mm��ʨ�yj�G�EGW���I	��<�[�V��Ⱡf�t�q�1�s.F�Q�P��Dr2ܴ���Ͷ����s�O5���C�M����7io�+O��#2���~���%rM����8Y=B�,V.,�U5F�I��n�i�k�Q\w�0*�F�'�T���XW�!ِ�5\v��B,30���O~&��ی鴌����JBw�D�BZ������<�!�_.YL�*o�9F����kՁ&��<���5s(��^QB�uL���Q��QTV�W��R��� ut�����ZЊ��(9��[����qS���b����r��S��ሒ���w�>��陥(����l�?9	��C ��� ��w��m5��5�����:����6� 罡���9��"��y��>a�n��� �Jf2##���R�۴���5�}���f���K���ʷR��$�} ��L���Aƈ
cd�G�t
�ʴ?�>K����D�b|�fʑ3�[�����A8�	�NJ�� ^�&P��@ZB�l!�*gJQ�`DM PVɏ�����1��Ҧ��їnሷM�E��b��MiwK����[Dw~�FZ��V��뤢\�<s}���,k0��"���)�������.X��m�t�ܗp�_�?{|�����*�G͢�^����9>	��y�Q2��&=�y���;�M���Ba��L��^��d�`,a-�v��ߴ�o�@�:�,��t�����Fs�= �	`k��������'��8�n<l��jd���
R9��7��KpblȰ]���αbY��~���k�k$)�!��CL&=�����V�ƍg�*ݕ~Q����!g���2��������)JIf[�e�{;&���qBQd�`��C��$�̊w��[Ϟ�'�!"L�[	��'_>̈́6�:{�ZrKPE�@t*N�̋�	�������D�8s�2�)@�p��82�u��y<�N
27Gԕ
8[Ĥ���4��0�P���i��@W�2�8��AS���I�lB�]/��tK���7�t�-N&�l�h�ò4�d�.;�2r=Wî�®��ů�n@�����Rw�>j�05��Vp��x���};vp�W��^RM��`)b��tr�W�'�� .�R�]LT$1��1��Y㼥Z�fw�04R�r�d���9��~�v�n�e1���#Yw�Q%�?��TH�ɭV9�f�ZӁ���*1�tl��'���8:���a][��FY��J/��׼.���*Z�^��4%���T��#q���Gi*�H��ľۃɋ���t��|���N�R6ccå�Y�:��蓚<تN�K'f�D����54�� u�m1��m�p������AZ-���ow�o��C��\iWl۶�g��$4~�-7��λ�1K��*�t���!jP�7���.���F�O�&8�Q��S/4x�=�Yz?�f�G"z�/"+�ȕ�$�qK��K�J��@} �H������f�4E���DU����rT!j�ޛ)	��[6�p�=���[K)�O����i�	�#b�5��Ku"�.*����J.Q�ermT.�W�_�*$"���5Ά�{{�A0kc�'W����M!�� o�*tۼ�ѓ/6����*��TV�>]9�