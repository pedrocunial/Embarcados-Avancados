��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cЌE���M ֫m��hE@P07�]���E�z�v�2B/�D�	��M�/ R[�G��,��)��^ނ����ۻ��z��j�W5���#�O���P]����_��'nW5�u r$���u����Q_��� ]�H�e�t���ڒe�I�U5����8X
�0����}����¼�C`$��pϥ�0�������s梮��J�(yi�O3�`��1���y�C����=Z�¸��$[ 8� D?+��*�����kT��leT.%�"���S���y� ˯0��/�Ӽ��Bv�8V��F����~�fMn�'�^.�q�a����;�ǫ��(zi/=4\���s}r-���}�wQ���Q�.}�\�1b��z�C�V1����P�*jZa���ڸ_)	f2��ݙK|9�]>��?�-SR�<�ѻ����`�Lzy�N���~��$J&.c�� H~0\��W(n��{�n�
ʤW���]C�����αe�M�o����ބ�l��������j&����(_ �wU�y�����R���)���e�蒏ڏ8E$#\�ێOI?�SɁ�<6���iD*�֦M��ܺ.ehAyƿ�5B۩6_~��{�B�O���%,0��Y�6~�-Իw���3x�Q 8�l�Ĩ��(]�Ԏ���	�F׺���'|<u�����P����֋�v� ;�>�;��� [+^��Yi�2�ݿ�`g� ڰǖ&j��ņ����w`s ��=Ցs�U�a>;��7#2R���2�	!`HR(��E�1&�p�%EmB##�j�J^u�?�c��u�$�ȍJ��^����{�7r�ܛȘ���u����
N��>�`�Ši���pՉ�R�I[����M#���M��%����p�5��)b	�p�tC��Av�N�s>��8��OhLPtLU��'���j�&b��㲭lW'�Ǳ[�-���9�P�z6��~��}�z�SbP��|l���yZ�!zǼ���^��?3vay���%�S��x#���DUM���n��Z��~GǢZU�N�118��W�z�VƮ:&��B�kt��v��m?<��� BƧG|����$�}q%
ʬ���=���Jj�z.<�)}�� T@� �����S;6�RA�<����~��%�7��B/�e"�1�����R����`ֶC<<X[���J�c�~�Q�U�5G�y�����