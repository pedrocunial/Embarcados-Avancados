��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cЌE���MuW�H��I�EyJg�w��L�Ħ��I����֮vt���\�Ͽ�ܝ���`A�e���`�c�m��t�õ�nq^���I��a�(H�V�F�'��7�;TugP����ԝ@����F�s�M�����P��
���j�;�����J�cv:�{�6��5��)����s�Ƅ#���6����O�_�M��O�gէ8�@�5$���(��tu���$Tv�lƳ��D[��!ظ�`�rIE�@���]x"N�C��W�*q�}J��۔P7 ��a�˩�W���ݨzq�Q�y�`��<�J7b�1;�[��!�!��QCŴz��JJ<���)��'�q�^�j�]�>�9��WͻZ+Ea4m�]0�7s����ɬ7;y�A���"\iL���>�s�p��<p.Y�3.]|L�5�pe�}Uz �(5�M�ۍ��MS�&.����+�OF}�^'�/x(���-Z��.�(w��#�S�@�)x44Ņ?���(�!��g�X^��|c�u}U!r'����=s�X��J�jcp>�S�b��~߹�b� �<�#Da*��m{o'�����l��T�.�RB��p�t-����`	���(�P;A|AV@0�lu`��jb"$�\ ��ێ������;.�]���:ۊ��y~\fɵ�IY���	R�Ov��Z�J���u��h$�+�
�9�_�)�VjY~5�!��6�ZnX���b){cӜE��ᾅ)�K��o��db{�c�34W�)Τ�6�GNa	� �8�+o/ 8��,�jV���#&�%�=��0��ɧ�P��f�IXi#���K=g� .�����'D+�c�;m� |��,�]-p�&����$�U�
�zV6oF�(e
���Hdq��ʞ�l@�S�*��	z��X{�NE�P],1��j�ݝ@���Rd��Mn�Q������ Y��bg�� ��<T��>y����9pf~z6��9Ēֿɥ�E4���󐩢�D��@�Z���z����6�-���]8y�RQ��>����F;W�S�d��3�3]v��S����!�g�.UB�+&	��]�*�;�#2���ڒ�Dg�l'4R��	�7�^�唨�^d=�Ys�$ؔ59�?[2]���</a�g��U�獬	۴]�5���1�_ʯ�O����p�Lx�<��Kȝ��rk���R'Cw�
:D��=� v-��	��]��*ĩ���}�d�wٶԿ[@�x�̼J����;��I}V��y-�1ɑ/yB��y)V_�v���g��B�������Rp��[�l�\�����-�6��T�W>����f�M��4��ܸLi6,�p� ��U_�M(j�xd��x�;�C�x�W'wR>V�h����J�5��yɉnQƐO�?����z}�ռ��Nӿ=U��[��4��˳�f�F�~����z���PO���p��׵��7Fb�jH��F���,k�����X�ڊn����oƻ��l֛�V$ܲ�%�'�:�.��f�r��XZfy�:�|�*=�7p��_v^6"޲��Ei<��ڞ�/�|��(��*��>
_7���vߐ5��=�b50��S��@M�sY>���75`�C�qW�)����C�Y���u�C~���(��տc �Q�pY�r����A2�z'D������:�:,e�!㫚;Mf�#��co@c���k��5�v*l�B���,����z�8q�T+;ujb��ʌ��G��6�}�Z=�oTx����j������2nQ-��W������Z�&y�MɁ��T!п,�-(%��-��%:�~^P�s�G�*V�k�5���3���X�%���ZE�U�m��҃��9iȤț��(j�����S|�o��ߔų��T���
��NE�^��v��|#�+���M-u��g��r�@5lP�M�6A��z�v�ۙ���"9#����zHt�%��Q���u�)���.�2����*�X�o�L^��g�(��]���#jG�V.d00tk�F�&�J�H�ʔ}�G*���w/�SѬ֍?�3�}����w��x#��a�=��w��Q�ʩ������ 0c�H]�7G��ˠm$iB���	��S�A毯����U��-y��o�FŢb+��V�o����疃�O1+��*'HȤ���lA9E��TZݼ'e�ϣB?�L��
������߅.l�V�	]�]���PT�ǧʳ�4E�|A�Ϣ�Z~����CQB @R��O(���O۽���w��A�~��6�t�^���}�,ϐWg��7�Ŋ3������U����r�}���"���˺�Tx逾i<3O~8%;8g�;yE{Ct�ҁw0��o��Y�a�?���|��Lcc&�����m���;�8��⏯��Ψ�hɡ{Af�IbČU�]���9	��	>����K�{���(v�#�uϱ&�ϕ�M�"	cko�g:�U����&�p=.�Z+�1��?��j=S�1	�5���.�Yg��B�K��B��f�14~P����o+���/H�C����y�0+��H�Ƅ�Z 2��ցV����t�rz�0R�G�L:]�
�7��f��i���� ��<�)5/4�@S�L�aA�w�J��P�f;Y2wÝ�fL2�-m�߹�?2���������j���mx6�G��(9�s��g E������R�uf�)����}��ky�A	�>�Q>W/Z��H�����V�g�}�)'��&���*�e�������ؓ�&K�ԴO�����?�;�.������S��*�<[��Fš�i�#�{�p�ќ#�ñ@��_��S�L��T���3���+��<�?�t�Z�5rV���(�TW@�['�}v �\���X��k�Ձ�r}��7(��Uʌg����L,�N����(�5]P���V�3��q`�-2r�vW�xL��\�?���~�թ�}��/x_�o�7�O�x����X+� `�,��z.�=| �����;6lO"z�{���Ne����׺9>e�J��,�N�z�|h���qm��qim����~�@�v���;p�KD.6<�t�~F�Ϗ�~aR�M���U<���b۟%Kаފ~b
���ed��EȾ�?�20R��~�ױ|_wg�������j�́���b��*KHgu�O3�U���� ��sj�P�;'LB2��^�%mGx"A��?4�N�Ӎx�c\�̯�:ս��ISB�n�6ꊅ�4��V�
�5l�)�i-���Sw�W��5������%P��.(J���Oy��0�[��b�k�NI����}��P�J�{=%%�4�'@v5�;�����x�#d�P0t��kZt���bm�[@�R$f��2����=���kN�(Fw�Y�Tԍ���ሓ��,��:��@��w:�q��=[O�ӣ.��Aχ��!�^cL�Lv:F�	��R8z��v]Wyh�_F̛Њg���״ƅO����g��c��������-���h��ڮdl�6��<�!��Gk�s#BB 6ub"r0Ɔ�Ѱ�q*�~:�2���� ^�QE���T$񴹥� K6��+񡓹��(��G�FۛR �|v.��f�G*��,��Y<��u�lSdW^�v�xQs3�}��2�P��P��ǻ;�5q�z�����0�a��ɿ"�Hn:6RB�ؚ�����[�;][�U�[��-�1�W9X�:�u����k�/�|�K��9P�n�2%�o焨����j�{!֭v�u=�.3x�/��ݸV��4����xT];���^!�,��(�(�gT܈��ϟ�ra�����������:@�Dɳ��349�XҶ���h��}vs+*]>C�����O̯� ;���(1���XF|~k�J9�^�-��d7:�N�U���Erj ::aM���4����r)�e� xҥ�w�U[�����ӄ��z��]��хU��ǅ�_�F~��d�^�[��.��h��Q���絣^�ns����<�.� `E������(b�E /�΁��Q��6��� @�wz���S/4��_w�(�կw]W�
���@�+�Iƒ�<w���b����@�=������xv���0A��ƺ�4Y��6�d��|c�i��	�h&�La/�����W��Jk
��f�h|�$�[熮�s�y:t�H��ݔI##��.��[=O��a�<t`ECv�@g��� i�7#ABlX�.��у��ϝX|���y�1��[��qqP�@y�w�@3������m���iU�]N���1����}��9����E������Q��m�������{��g��s�SGj2���B&&��&��n%W�ґ��<͕�D9�ߥ���#����O����>�j�#J���5Ĉ��u�a5t%,-r#�>�߾B��D7<`��C���2����/n��dV\.k��a�aUt}����Z�݌��@�L�zx��py�گ2���9�t�;�c0� �u*A���;�p�T�K_E��A�<�AKp�Q�����X��
E�oUƏ
�����K �8�;γ5��.���Ar(��sK�P�f�Q[z/�W�׿���ܸ-����w���ufD;qi:�N<����Ň�fd���o�}�Uc�
OB�
z"���>�}C��Ăf�C�寄9��L��o���+�Oc\ 'q��;�ٯ�w#�P�Iv"H��P���T$�3� U^z��A�����xo�#��7Žw�zWt�Q*A,�-�eh9�B��k��(Xs����k��V��0��Nj4%ຽ�;�ڥ�*�¶�%:!a�����!9�Z1]��\���/m���k�;���Zc�o�Iv����9-�ե8B��3�0�BEю=�&kϦG���x���l��k��_x����F���v�`�������;-��7��+���n]=�ʈ�sio^�kA��L�gLvN��UY�Ҩ~ui{F���}5�K���Q��Z�?[�bB�Nqh�8���ll=�,��P���.�QX��"8Ɗ��0���߲	�+#2��B|"��	(���^zP�B7��`Ӽ?U X���/���D	>���F�,�2
 ��f���������b��fLލ�?��̆ƒ՜*b��b!W�Ȑ8�KavW�drJ�d{Y��֨_NI�M�*o�V���L��u�L|*_R�?�&@�V�貨�0�#��<�\J��b�&�~)��^�p�ƥ����9A�T�pV�V�tJ��d$��x��� W��$��[c�1!�g۴aOxe`^g���z��S\��O*"/����MP�=	�Ȟ�e�8h xEZt�AZ���hP����w�
��dx����M�bb����nӿ��կP6=`å��!�\���7�邈�`��L�Kz�VS�*�=)b�֑���|�*Ep��o����/���H��l�+�}�e3#o�p?i���=Hք0��[T�������a�����\�Ɩ�bi���
-2{�TI����f�00eQ�{LE� V��&�`3l勑05�M��������RC
���-�|��	�0�R��H"�
����e�a�����\�)�,���Ŗ�à0�s,��Y�Ԡ����=�*���� f�ԅ�;�m�@����N����;�5�xK�Pٍ�m6xٰ��<�Y=��ET�F[���R�y6X��*=�SK���zaY��V��@8g=C@�y�D�Gv4��s����asUԽ+�_ 4q�����SWQ�tMwM�������<���WH> ː:����IQ�(+�S]d�Pw�G6�ř�ľ�h7��Lh��-9E���� d��P���͏�$yL|k{��Б~�,��ы�?��\��cvJ�9S�SAoY$B%TO��ɫh��q�0L�T�s�u3�]���.�B�]�. �t��`��r'��T�U ,v�����x*�m�x�YN1Ao5"z��ٙ���- �xX�7:�%�|<�aɣ=t��#o]凊�bU�l���{	&:0e��2�Q�誾j���v�J��Pw����u6��Z�p�����Sj���1��Q� ,v�,�YK/oh��H��yq,�<�Yϋ�_X��}P�c�⳽\a�t?�\wdĻ�������-�b�F�]��qg�"� a3��5�l�/��|{jO�u�� �̌����g�g�in���6h�Q���ܑ��Z),"�M�W#�(��Oq+ �iM6�f���C-v�r�]�F�R���������"`uC��[QN
)�{�*��E��G�y�i�@���[��� }��*	����9�3����� ��/��"3��M�鈗?�qjt,K���~��){��}!ؚ���@��N&�ODx����1U����S��6��ǹ�A�h�>��D4 ���dx	��ߏ�3|�z l6q�R�{�&�;�=9���C�F7�����lTҟ֝i�>����yA�E<�>����𱡅�q'ior.=ZN,<�0O�8*�D���!:�TDԘ|)�'s������̲-nu��1n��o^��l&���Bf�}��N<GM�	���]�1>a���D[�:��gr�1ݾ�s���2�����Y�� hRnE+<���㊢r�Jz�!=���X��OG͢�0	�/7�g:�US���2^?,�ߪR��w�J��"x�io�-x��O�<s���� B�y��s���������o�8���	k�����=���"��χ~zs���#xA(�D�W�V���c�XR��:>��K:V����jvZ��x�Y}���AB���,uZ)�d�끍c`��.垱�/����5ݭ��w|�O��R����t_�1�y�a_wxw���,���u��"gHخQ�-DU���\��	)�k޳?z̒��f-;lB�h{+3o�(�P����;!���4��E�x�-���eV��$k��P ��`�}-U�h��O��7:dT��J����[��SΠ�H��*�EH�����<	.�%�G4U�K9_��N�ބ]��&��k��o�[�E��Yq˷*Z@In?vW���Cfmu"3L�,އ��2��[�жvr����qY�9��u� �+�Պ����$��j�0��. �ё��L"�_�"�ZǈN���oO�0�+j�V���4�sY�>ɥ�E<Y������S�yTq�Q ��c��,�pL�ul~eA����bvh���jX�����-�;�޳%`3N�o�s���c՛u��x�S�6�G_dX�qw.{G�l!�9v�H?*��z� ������%�G��l��$ڵ�`j�*I�k�%2����V^��T��j3Δ�o�QԘ�.mQ�a�X�G��~�K6�7����-O���n5������b�_��%D(D5/�&�us[B#G���J!u)�Ui|��)�� n A�]$���S�G�+Ά	��hQ����d�ѡ��5��T��ဃs��-�C���QK��y򛼋Mz��'[�-�D2�s��H���^�%��i��ƃ��ە�4	�X�|�[��6��j���LƯ=p��p:$�����
��a�D��1�L�d�2'H�(b��:�E�-'��Ʀ9����P����hܩ�;�`;��������lm�i���8J��'�)Aw���~�A{r�Ie��ߖ���ʌ>�r5��͞\�_Fkf���̣��ćB~Rv]c*k�A������;����%��ڈ"��nR��bʆ%�h�ke2�l�ޛ.��1{��E(	��)�1�����XF�P����$�3�4^���j%E����>!]��@(1#�%�Fa�CNԢ�q�e9�������k6���� ������/ib�+����Q�%h�?96l$�b Ǚ��#�D��b��h��LO���"/i���-���)I��Ɲb��D��1�	�/k�M#n�V�0q�VC�jO)m�Kv��r�NH0�g�'zݟ��9�v�%�ZI��@�r^�yLL7w��/�Q���\����~��م��WG�`	)�������>y��)���9ݎ�=�sa���կ7�!�T~���U���N�X�!����_Y 0S����@�r�t'��ݮ����Ҩ�����ݸ�M���+x���~��`L�/�)��A怤X���q������+Q�W���X��9v���K~�L8֔����,$y�L�;zY`��,@�V�!��t���*��C��@�1����̫�E�6���=h�PЈ�6>XU�p�����9��%(�L
�:�>Af�Z]�]b��;�q���z�������7 ����Կ��i�_�<S�w�����oց]�s6�6����K�sC�q�H���й�'G-�ّ*�6_���O}�%���$�#z��a��0���]*��\�O���\�ۏ���}H�Φ=&�8W$�J�?u2]4s2�jR��p�;�q�A��Q�&�� �BRN�c���XH-�X����%��\Ἰ9g�����-�ٳB8���E�ˈpZ�}n����T͎�A2�P�ܧl2&�E�g½p��Z�d�+�kw*q��s��	�	y�#�{�qTl�N�xX����I�b�b��<�ow&ߦ[Z X�����탡A�X������3�����/se��6�,�Z�L��R��+˦�M&���ըBR�I�)���qE"I�-���(��XZ�a�A~�u	V��l����ʬ$6����wA�UϫM���q��w0ɟt}�6�}��z��ݷ)#9K9V����g�T�w{���d���}Q0Ӣ�4�-��{e�c�L%�o�o��7����3s�l�Wix��v��ٔ���O�!W��3��Q��,����)���Ēc��Mgu�hG�&z2),�Xjg.po�,7�E�f�����P0�=6Os_NR�45���m��Q+���X��3s�Cr���f��Tc>�(>Ī���_l�$�^�uly��P���Ϩm����&�s��F�����O���[���7v�\�"/�U�� ���o�#E0�O!,f��Ĺtsz*T*�.9�a�lR��q���0kuf�`=BGɏ�ʲ�ͷ��+�?���A�1X�|�z��mj�(N����+���a�+���Yl�C�k���䒾�L�F��w����D~��)�� �4��w"-t�M�j�<�`T6��S������]�K:����}��0�e�:��:Ce���m�V��}~���~���}{�g��0�7�\����SVU���Q�Μ��]L/Lk�*�X-����~�9��\�T�ZfO>8)�]�����ڛ�-�e���X��r�e2zˠ����Ψ��Id�r�U'K�I��������A��b��)7ceƌ��4c��|�>��T��n����՗��0γ)���ܑR.�9ûfx1}���Is�k"W֊ٞ�$o�Cn��C7p��S[���6�+~�[��n��t�:��)Z�~������u�o!M���أc4��3��E�8����_-o5�$@τ!&��J2,�,���1�� )�(���<\�ޖ�A"�O^�9.���gi`��}m�}�U~��dK1� �n���*��#���K�"tȕ�f=�ٹhJ�3��qγ�qvC\��am�t�
K���)��$���E�D�=�O�I��/6�	X����?S�ץ�/�1Y߀�#xn�
�(n��5�״^��h�8�H�����o+?@��Ƥs��>�Xg+��Cqw����-N���d�M�&E(�z���s�!I�%K4�	���T�,�L�M�\���P�u��CQ��L2��b�j��x�?���3���������~����P��a�qa��UP&R�l �F�u�xT6��� y�a|�A�Y��,o�WR��Jxa��]ՁQ�OIN8��h��=&��7�8����v&� �0��	X9��f���,L����~C����LR
{˔w���D���]�$��U�;ć2*y8kuK�AI�ƴ �ڈpZ�[�}��)��>$X�T�� �����ʝ��.�6�S:jHa�x.�V��z�RP�|1e��U�)l�=牗�YɠGP&�����X)�㬹�j%���t��KE�~�Ws4�<�l1z���ؚX�M^ü��߽�P�J|������csj!����'r�O�����8�uN�H�xo�u���Zۍ�U[���$Q��Ҷ��&�B����c�7uFS���9Ǆ��3AP,�k��DGJ�N��+8R�Ø:��w����Y��ħ$��ɛ�+����Dq2k|E8bE�E�=����lwۅ^��[{gɊ��z���^�X�����.�s����;�~�+"��+0>��`���R<[䪛������ [{ ˫��a���w���n\��pJ�C������
H��8���'��KΦ;�`�3k�}����-�N����x&��R�5�Ď�1���m$_*�7�`�~4�i> ��NYN1cwK�1]����EڜNH��b<+o�Q��-t�T�� �C���y5R'��m�º9�5mq�Ջ�YQ+l�[��3,g�Á�bP�����+���N;Vlx�S'��� ��@V
�G����|���4�RC��1����XuN�0�G���w�'��C��mhv�r�Z�@7�B�Z�w�F�D\�VGP�k�n��a�i]��P��KuS��^�����=�@�X
�&>�%·�L�Rn�t�υ�"�:G�H�������gN����'�l�A@��$��(N�e�	�B�_�W;��?_�vyWMA�a�١+��i
 �M�p�HJ��cG��1�ޓVI����:����Z������6O�q��d��&�{�x㐊2�f�Bm��h:�UӺ,��ZXޜS���?Ļz�ZO�Sk{Z�c��࠴p�YGƒ���r��0��s� x�p����ړ���6��u�ᛏr��$(C����^Q��4�����@nFD���Q�X�?/q��yqgcڮ�����$�y�m��D�(T��߲r��{����%����
*$�+�s���l@�Ox�*��rz���׊��nWI7`���M(�`HaÌl:}s=���U���th�:�?� �s���W�f�xi
Zs���ӽ��G{�1��E���(0-���>>�l^D,D����`M�X��}m�Q#9������߃Ia���*,��"=D@Q�"�l�	�Dڢ\٣�!O���b�g,�,iP��n�԰t�kǌ�W�ȤO4Ɇ������fxd4���?�m���j�^�L1ֲ�;m�Gwe�r﫲��}[(4}_f%� ��;3{�(�8��D,�x;&��kD�[=.����7�<)!�&N��h�R�ux�6ĬNbq�+�'�31�M�;�wn�1�v��͐k�������J_*kٮ[) sD�k)!I�^�©N1���o����=�s�ƶ�~`Ʃ����A�7@/���T�^���Q7���!�~��`'#�_bar=����}ze����*t�V;Xձ�-���_N�<MN3IBKI}@�e\Yb�v�,���>���{�a���h�CWꖘO�$�5

�"  xOd$�6�
̝� ��q3#��/w�}����x�~��<���e^?��e-�J��XJ�����AM$$c�$̌R�e����F#@(J�q'��4���W%�?F���lH��8k[7��+�<Uˎ�Q������ x�Ԛ��SL��s�@?p��čD[�TU|r��?�OI�R�+b�,����6���"�#xv���"�}f$Ў.�'^bt�Q˜������Β�t^ �aIub'��r����xJQ�{p�9$��<o�5|��i�����x�l��P<���Rۓ�z1/d�gAi�"UI� ���\�:̸qm!�Z[�@O��3����\���Z�f� {�!���G�i�pb9e�2&��x����%�y_��C��49,V�n�<��y����l{�F�w��
��2�R���Q��^��}��Op3�'�@Q���Ƌ��d"���7�1��]�ě"�`��=��5��p<%�k0 ^�*��#��<�����[G���󏞮^��L*p5���y鎻�s�J�>����F!o��� ��fŇ�<�EG~��D��D�ٚYՠO.��D��|]�auኘ���uȬ��$�3@�H�|.�����&X�qDY�~�DI7 `��y�V��	��Xk���]Jv�<�}�E�3�؊c�m��B0�vö�1���%{�fF�(��J�שnM_�կSJy!�DUAq����o�|�*�m9�E�gm��5X�j��):Q�c"`���}�����%�%��W}�vw�^\������t�;�V���`-��$d���
7�PPk�]����z���q-��m��f/�a�@�j|��P<{!-�Р�oSyN��p���^P����b��No�}t�=�;J�s��g��"4�lf�k�oӃaY�*��A�8�Y(�!n����Zw� 8��(Ǫ����UI��WW5
�,|ת[��b�ݔO�Tӕ��`���A6���4�JE����8Ij	X.��:7�a�"�Ǐ�G^E+�rSC��S (D�+VE��aohJ�3K1�+K�!����I^=�>m��-"hZ��	�N���+���uo��[<�����~O
z�������zȪ?.�Zp�uM+@�*y+�ʲ=Amm" 3���!?�y��C�$@�j`|�kB���Y�Uq�]h������bg���=����}��sL0��ٱ�̌��'��S\�aW�Ɠ7�hs�V\�=\8>4�ā
���os2�ԏ�����J�D,p��.�<��z��F΢h��(��)����B	@8��
��v�9�)�J7�1%K--ҙ�ԣ�3֪�h�bV^ ��;�]�Ϋ] ��q}�-�[QvP���y˷���h�&���t���r��2�?��#��
����Ԃ,ϒY�{�0#�h��ax\�^.T�u yN��ւ�C򤸏�!��Z�	Pڽ���������ձ�.QD��	��G]&���$o���׻W���Kn�(j�y{gըSci�������0@�3�d����2�����Ou�~�.;���ኝ��lQd�-ư�J|w�������_�9���X*�ǉ����}����%�ja
	%�W�k�	Xu F	R�X-c������6���h�"���3��,`0τkr^������M���K�n��Q
g�jRr�I�s�M�95�3��-��{�0F��1�ܺ���ƈ=H�Ƭq�ȥ�4��S@��\H���y�f�TW�kY8�j�%�D���?����a�Y0����%��u�=�NV�v%1]�����h���S9S�QZ�{x���W]R�$ܼ��:���҇��-A��^�v����^
�9�#ݎa�1iz�(�c�L����y���Na��-��~D�}e}hl�C������D��Sʋm�MB����c�\���k�+fM��p�:�\8�U�~ޔ�g�7侌p���)|���3��Q{����d�!sP�yG�%����T���� �ku[����=�]m�ՕJ�0�h1�߻��α��E߀�^���� �CU ��\y� nĪ�����e�����eCr�q�(Q���M��Ag���"O���*7wO��V��Q��O;M'�S%��5&��҂1�A����h�J�20��J�>s�S���oz���ż���/$���w�'�Ǐ�{T2�p��}c�s�#v�>	�u���>�ѐN�4��+�6�t+�z���B����Q#��M��s_�-b23K�/ea�K���eƿ�S{?��\r�˨�3F�F�.��^�� n���?�,�k�g�� ��?�5�hEi�9$��|uY��v�~��sd��HU�A�i�l(�ʁ���ըOS�Y�3��\��Z�.t��_�'������H�o%M��6E����W bK\CW�f�2�A-.��?��@�HVM�y1S�J��{?2�����h�S�7K��g���mw�&wx�3oQѸ�:�dp��b�,��Q _��1)����˿�ܜv��wl]�\���U.`����0�C���p}�*z��-w"nb3j��<�H���������6�k��$�h\�Tm��q���p�7<ee������X��0kCG~}����>$��e���ut�Ee{�2l�Z����N߹"�E<��bV��N͕a�m�����j�t�ڳ����f����Nyd>+#�X�V/EP������N5e���Ji�֥&/�	��[*�?�U�V-�hM.hKܓD�}�����չ({o��f��d=�b���!�Ÿ��}=��`j�\:1X[�+5\^0���%�&{���o�r���U�{q�Sc��|�t@Y�xJf~ʩ%D�P�C�A`��,�=�A���uhL��y�eΞ2���҅1�_J�1�E}��MJυ���׌�X��+�h#��Z�r/L�4S*׶'$�P����q��(�.����0��B�EJU�@��I=):�̲�A���K'#�����rpZ��a�y���	�� c�]���}�j��Zr1w
[�b3/򫸟�fiݰ�Stq!SBW���y8��(j��S���"L�Ua��t�B��͸('���)��5��K��Ȇb��9������4.@�ݨ�\��q��O�"���fܦ�	x�?���v��X��eq��#L�G
����I��X�$�~G�|L
ًY^3%Z�p)�����qJ{��X�!t��H���VR1�^~8y���)�u�&H����l�2?�U�x�Օ���������5��6LP�n�Ҭ�,nA����!�,��9I7\�Ga .�&���P����!���[R \��.��'��XuC�*�������*�A�7H�)�#,n�&������ެ�@d��n��ʂ�)�� Z�2��@����Yn�uc�(F������~���G������[�n�����/��\�E��A�`�ʗR��B����L���\��O~�,�	�5_�<M�Ee�$\���{�$`x۬�,N�����Ī;O��g�%����(��6+'M/a���",D�����*0_d�®,~�#~�1*�>d6.D
6z�ŤzGy�˙�:o�Wo�^�]F������n�#K�5u9�_oE�8��(����RV�ۀ;3�$Xyp�g���{�W�
'�%{��9%,畹~�l�˸j] �6YsdzĪ�h9�����T~��џH����i���u���5<kT�a^]��83R�R�5��R���d�c��JA�q�:%�X��-���E�QL���%�{\f�DC�^�,���ÛH��Q(>~+��o�1���]�#;Ȳ�3
�c�Z�q|ů���Y(T��Zy��C[�E@������S����b��`��rx(6�[W�Z �}#���<\q= �|z濪������ 4 R�P'�ƆlP�U��V�ӻ���pb���T̬����ae�>��y_�t����Wx MbY[	'Gu��W$1 ���r��:������n�v�(��&zS@9Og"�:׮g1�7�h��#�U��P�2o(F��!���&��f��[u8�m�ꌾ����a:v��|or�3t���ۑ�@O��f 	6� mSW@��4����(�lG�5�P�
�ŕ
�ژ� ��o��p-b������!]�U�x�A�ِ�;�b&S)Ғj�����	8�s3ֺ�:���mƠ�؟7σ�ד���#HQH�\�f>�_+��]أ��۸��ש��x}�0�λ}r'�S}��J~�����[�o���w%%{u���Q��c�j�JK[���A�wѬ��Q|�:����#�����&خ�I�x��_��GLx8!�cr�J!��U��^�%]�1S��~�4gt��;&��F����<�jGR�r���i�&1�k*}�(��_6'�Տ_DhL��\�Lq2f�ڧ�� ���q�=Y���K�,�kج�t{���c�������ec@����𪇳�8x�w�2ZV2O��~�5(������O��"�v��o&=��v�k��J�Ȩ��~Э	۳�J]�j�->���0��4�+$.�XR3q����ah��Ƥ��ܪ��;Uz�b��.���!$:�֠P �^8�Q���*�Ve~����V� h2�{"�P;xI������`~��o�G3��U
�l��A+����B�"��H�>O?��f�U/�N����X�O���
��}�I�����D	H�f����f>�g�a���d��np��8Dwt��	W���wt�ym�dS-B FX�q��_/�vzZ3���
����>H��Gt������ɩu��������z&�����NZ�`/e��b#���Jm$��NXJ�����Zcwe�Os ��z���i����v�'�����T)��}��c��j�rQ6��S��䟺��ә�(��I]����������3���	sO�!Ǵ�Q����а��1ja֖�[X�R�~�7}�v�C�������7JJ���i�T�i�*G�?1�� my�K�"��3�h/w��Rʄ�����瀝Z��<K��f0ňx�Y��?z�M=fN�&c��䣨��m��>��'Oq���d+U����� ��Ӣs"�ٛ#��n���{�JWx��4gK�����I7ٚA���G@�eK@�T���_E��P�����5�$�\RXL0�7B�S�dn���j���3��Й�K�Ǭd����Ɋ�A�/����(�*�?j��Y䍨:�bV#�Rt���H�8�����AEG��-�S*ޢ:[��38����r	E������Ҷ��X�J<`��R��C �z��9)� �hHdf��	ߥT~x�J?����o��,���Z6���
��ڔT3������`�'0Ju���F�ǯ����n�sf�ߪ���7�%ȳn���)%Һ�[�!z�k���� L����N>��Kf\)N��mO�]2۰�p�`�V�W�3�v��~+���ȋo�:$=��Onx��Jb�O���Uِ)����"�jiǣ���١t��dn1J�n��~�?���Ny�U��k$Z�z���Gt���X�*�A,S$�����\�WRc�	��S[�q�Lkh|3�%�y}_�%��~�0�hnlp4�&�l�x��撰W[�g�(Bh�+��z���vøh)ś�@	+�R��
f�A�	ѷ,��Cބ쳛�����伯E�_d�p�d�?jt�Y��IV�o�@
{����T�|��,�r�%��y]��F�Z�����<��ɘg����
�s���[���k�[��`*U�x��`��5���Ϻ�3��v��}�N.�L��+_��jPM�̜�����ږ�%#���3����[�t�dX%�l��ݏ��,�ylOs;#�r'D�y~�I�,QTi9%L�}V��9s(��U�Ti�M�r9_���Rl$5��ጝ8���?�#bo/��~�!Ɏ2	hk�$������eq��
�����8+��ۨ�x��d���yŞ�	��6��*�RC�c��2٬��r�ʦ��R�l��I@4c3s4��[Z���3�to⽩��h�b��z��$v�b7���@GH�U½����ܥWr
�Sͻet��бcc�q�ׄ��\�ؓ�����5{㱙��i�n�Ye5�-)B9�	��[-�7i���H@%|�r&1�l����(���k�Rͫ�z�����>�kF��S}T�?_�a<��u�L��vfLQ<��#��b�xs`�����Yq�������4��M�q8�q��������b�a�$���b��j�\�۾�iw�~q���`-zB����=�w@`F�{X����_YǄ�����P�	� ������ԇ�r}V4���V{�3�RVH&��2���������7���t�����p�vg�v#�;�ZӫM0%hR`N�E��hȫ{Bw�pĔ5D��5���Fِ7"���9�H
OHw�Djp�3��A�b��y��Bjvk�(l�KKD!qu"Ow`�h�~���T�e�5��drx�����h�@
��U�x�9�)/FBT����⊀dE�Nk��2˞K�I�s���QPq &���\���sy$2����aq��^�k+r(���L�L��%�}�6q*?<F�oK!S�
�ʔ���S'{���r��<����y[�w���GA׈��8�ŢB�s���m�ǳ��/�e��Ѓ������z�:Cr˾*�����=T>��?t3Ry������k�ه��h�cf\{F��LNp�zh���,���\i3D9D�~��<`�:%�=�ꥫ��|�/�)�؜^ʾr<�����	��3E����}��ā�޼x��a�j�ա�/��d��Ag�[�&����}�Ɋ1L�)��Y�[�$���1�t{�Ѥ�T}�u#�K���C�_��i"bT@�y���E����j���������If$yv#�)�O�.O[W��.#hb�V�C����7�SW�|�M8�[���)�.�����T����0l׼q�-��}ݕ;�B�hq��o�KOv)�`$T�%x5���j���O,�I���!�n�3�tb��ƔU�\ht�ePJ �CĶ6���%��9F�j�T5~�ɼ�נb�^�4� ����L@N�>��?]#Ε�f%��kw*�IFcV|�Z�j���J�UK�i'��iQV-��xǌ�̶�⬟bY�P��h,�[X�Ք�i�3,��y���Lv^^r�%�vu�>% b+����������e�a��AJ"N����R������@���� 'OEJ��b?�)U��-�10�1\-���N.D,X���Ӕ�e���v����M����a�E�Q�pN����<,��N�[����wvL�����iV~�8{���dڜ\���^�+�*k��� R��
��施��k
��.	�R���_����@[<���R*�ҍ����Q�] ��u�/��1��6�+2֞Z��_�z���Ln�D�a{��r�M�F��1P�C�al��o�D��.d��~i�>��Y��(B�+�������3��F	˕�*�t���d=��{��6CEW(散w�ǥ�6g����فw�w]���Ȟ0ڧ�-ie�	�7TxrҔ�X��f�,m6~�!�~�Ԭ��n��r�JC3S/��;
b�W6���S7&�!A�9x��������:�[�'_{�������$-.m�&�t/ +Ⱦ/U����C
�.Y��D��7�_�����g�u��uL
��
��٤W�1�ĕ����!��H$:` ������&$BTnb�S|J`��T�ѩ!��p��|�����=SkoZ
�	�}=�E�ۈ���kF���K�]�)!�r�hɭl��/��紏�J��̢g9c�Q�~�_�
2��$�}�{U/�6��u^J���iC߬N�y&ޖ���1X��l����i��o�=3�a�vCM�)`�ߌƀZ���.L�����Kh�2`��^��#6����}�[�6�E��A�v������[b��w"1��a��l��Ŵ��SM�4_����'��3������EԐ֭Z����ȵ���w\�g�zX$F�^$\`�m�&��RG�@�Q8ai5�{����~EMH���58�7��7F�e�P�I����|�2���W8�X�8����&����XV��O�-^�=��{"yT6���f�I2���Znű،��\�-/���bG,����7o��+�9�Yuܛ�@  �����[.LL��T�(6�ע}� ��Eő�3[���6
�z�@hj��3c\lCI<�o�1���k@��t�tal9d{E�X���KʮQ����C׶�=��F�I���3o�j�9y�ܲ'���`i��.e������'���~��C�P��ay87�QllwU������L�tw^&���!ɭ�d�����!6��(n5���Ī�����2�PY�ڹ��K�XU
�Gl�ݪ#����:s6f��mߋ��f�)�Kb�8��N��#������`��?��λ��M���Ob���m�n���a���o�~,"9�D|<�^��(�_Q@�������a�h��
�w�j�1_�.�p���t�?���|0��k\�u�g�5�WH�PX�et��!���#�e~L�g��BS`� �k�*s���q�T!�12��|/j�J<0DҊ����x9	>�
P���D�3(=�yd��P� �8$��/c�:�:Z�������^�P���1��	�o���R�8�;�L�-���Wuq�uCE;�`�NpQ�M�i�_(�A����l����JU��_r	�]`�,��y��S�~y�|������z@]CV���ٲn
��{�5�����H�o�_�c�fc)�#^x~�\*�O�b2���H�Mp]�Xz�v�ܜs�v��F��ܹ�0t��{M���p^e?�H�T�t����*�6�1���� ��K� /�t�@���F�B�����8м99LM7-�+������̓a�I�ϟ4��V(z8(��6)�G��л^7���q�!g2�����.�l��̔�h�b��4����y�+�͝ߖ�f�F^��5��{s��(45��а�6��>K�ZQu��Қ8�C�5��M|8�#+)c'�Q݀��^�w����->�Yn�dG	Po �����~��Q���Η\�7�,�����n��x��ո?���������*����;�{L{�#A�f#"E)�ϳ��)��^�9����!��!�"������2�
�����!�0�����ӭ�A^o����=M�������(A��֝�Uou�ةVT�zf*Z'����Ҫ�l�O�FV,��7-��A�([��e@�k}��ȣX�v��:��?4�z��wP�o�m�</��ܞz�R��XM���QE���'6��t߲x��� ���,[z�9��M��^5q;�y- 6�`0]e+�E����l��` �@�	ߢ�u�D���
+%M�<2�g�i���.J>=F��vU���g*���+��n�I٫B�4#|�@�J�w�]��ﵬM����w����	���y/<=3�w)�OG��Ъ�ҷ�v�4;�z��s�\�(v��wU�=�i�6�������Pq��S	����)���3)ġ�X�^�3<c�ڟ�A�������V�Ek���g>�Z�����*���>����Z���@u5e�^K�G��Pf�Y�V���.���]���1B+k[�exb��;TM,���͉�%�14��m(���ad�ٵ��\�|��3e�B�v\�Լ�3�Q��'(f���9�W~��L����bK)�cU G�=�ԏ
D8�
=�B�8H$�7�Q,*���CQ�����('��][�̹OP��.>�E�*&><CI∮�&X�-h������[8��F�����e6������`���T�܏�}"Шk��b� ��-nD(>S��ޯ�	W ֬\��*�>�m��};Be�L&;ɯ����ͺ�!@��������4�n`R�荂���B�#3?����[T����qڎdC�R��|z[����Y�&`�3�CS(��A۪�~R�e�5�&�@�C\樺��Y��+]��<�`X�Bņ�^<Z�šD'���Ѭ.����\�Z?��U��8>�� բ��s�ݫ@��\�j� =JP��$W�|E�P�o���k��T�:��\f�y���pau~GbQ,R����#�������iVI�ǐ2ƽO�O�6j���q'㙪9V��Nm#$0��� 8�ȭ@���x;��^�6�[���7�AˠX*�;��{2�|��M@Yp�1݉.^�*��ٲ'���\"JK�]1׼�3\�83�.�Pl�~��`�"�K��X���!��±���c�${���:�uQ0H�"�%"	1��t,�����d���7��s���5+�ǻ#&���uW���sEa3�R��ZY3�� 	G�����^PE�yp̈́�1y����k-�j��W$�i�:
I4Q�]�f�!�q+hi���^苦ʺj��<a���"��c;V�Tͺ�[IB.�{7]��C󝥴�m�+1�R��u>/z�ULA�q���v���6��x��l���p����@4,0�����Z΃�9�S�Jv`%o�
�^~��C+�����B�-�\[C�&�����hd#Y7��Z��&�%l�n!�0�
��]I1[<��L�œ��ﶫi;���b�X]�x/���u1���y�4�O=Mm���w�8�<n����@L$R����w"7p��)�����Ȇ�b�����5��}��`�/E�σe�a�Z���lzJ���G^�@���,�/����
�2�4}E����ǡ�dEIs��䈀�A�N��^�����	������Z����t��Љ�@��X�ь\�f��d��JvUd�L��/�c�L�i���TE��rq���6+�R�y�*b�w�4�Ͱ����'��g����G=�P	��4��S��c�}OJ�x^ǇH�]leT�y��q��pL�J�TH�<���#V	����F.�dk;��ϭ��l�) �����`����v����K�ۘy�u6�&iS1�Z75a��o����� ���<>zh�����31UaTq�M��]s����T�:1�3��]�b9.����ň� aR���7P�`�Q����3&�?�G�\-��z��\6fK'�Uˑ@2y܆ �߽��!�s�w��d������@��ˬ��i"uЌ�H���S���6F{k�.!���E5��~�~����q�p�V�������z�G)�p�/�v��	Zc8?�z�s�vw���q�[�a'�a���BB����Z�"��o
�p��}>F�Ih:�𢇱s6 �oT1����%����)	{���`떳=م�U�������1��b{)O�<�{6/����"�_i ���Zۏg�.��iˠ!��Ov�H�T-�I�H�#[(>��6�����q�b����N2�<R��'ix3|�JnX����_�n�1+��;�Etwe��V��;�,1���nJ�FlaΑ�V5��C� �Y�O�X!�i��H>s�S��<��aa�b[�Ўr��>m|�mx3	�(����Ҷ�F ���⎦���0~ +�����/r,$1:�����+�6b�������G�Oqc.�]�̋�r�--D��M��Pa]�E��*�g+�b1�L�Cވ΢��8�Ï�,53��nu���@2 ����0��u)������w�p2�D�ԑ����
�[�\�Ǜ-+�v��t��@9<�0��C�J����l�`�T��[){GB\�����ֻIT���mDD�o<{*���%����^H�(��ͭ���<3�K�����ʄ��ݴ�x�C�},12ѯ�(�I�^�A�`T|���4}�`id#}���.Y`l�o0��s#��(vƓ��XϤ�"�P� a٤�����\k��f�T�����2B-S^V>�|�����(`j��ǒ��ݤ�KR���/<s�=%�B4I�$8�5Ȍ���/.�ء�Xg|����"+�����lt�����]��ls���9�5nH fKd:�*�)v��?���	qS��1���A��4�_S�'�2ޮ��+O�J&��q�.}�3�aܚ�z%j�y�x&sT铃�j��d�n H���-%��M+�|�V�3���0����m�s�w�+��K�3��i(�	�z!�j���l"�ۢsg�-�c9��&Լ�oآy��R ��ߡ���l��+_Cʫo$�0�G�mĢJ�j�h�ݙ:#���ߕ$d��90i��]��k��q�9o������%����,�n�ө���+]
R{�4X��Y滨�O3�y\^8�?:D�an�r2�d�Y��]�M� ����k�!W��'�D�9����={�x�]�R1�C@�����;�����*�i���C���~�JR	��4�Eh}��L]�V�g��En��`��R��I�JZ���X��O|X!P_�g;�W��4�ᵤI��_-!��yL� q�C-�V+�[(����E�o|N�;__I�֝�S�>J�]��Uߚ���֐��@�B�#XZ	�a�z�<>1��
�]��=���qW����R2y9R�\��i�w��Ī7�Ւ��'�ʓ����T���Y�t��Y�o*L}(_?;�
����R��r�2
G��j�D�ON#��'�%��$�l�[��"�ȩ��W؄ֳ��/�W3,��I�n�%�"L�%�ϕj".��Qo���o>=��0h������o�p�4;�[oD�-�� nVL���u��e�� �Mf4ޖ�4׉����?ɂ̋�O��1g�KI��O|��.P���y��H$fY��ť���#�ǈ~�n�W�T;��矘^����/̌�FNt�t!��3���m�}.c$��F=���7����V�؏��>�VgE�e�z�!f#�~�dmt�ė��6B���q��j;X9�e��u-+����2p�W#��;>�����Z�T�4�N��2�R�Q!G$X�7g�\So�UQ�����vYnĈb�Wm֦yR�d�J���3sl�؍ܩ-S .ޠ��d ��A{��Ƹ.�5�{Lo+��������ǋh�+�X��4K���m�M���@���(5�D����ous�����}7�ٲ'a�)�:�:s�v�.ǹI�j���08�
��=�r~@�Hf(�g�J�:�/� x�-�E�"��9�j��#(�b5d�:6�.�uF�,��U7S���]�tk�"y��t9�uz-b�g����U��3�+�dc��"N�X�*q�"a�ϗ���)jل� ��e�Y�6 �����Z�X�k(�4��E�3r����Q�u�A����oA)su���;���������x���,B����;0�B��|���2؇�:�G���%JQ%��.��k	@�R����֩�;Wcp�����I 6��αL=q�A�0C#�gU��Bȳ���&)֝��b򫎓&>%�ܡ�P��1�c2�>B�D�XX�,-��qi�Ut<
X�5�߂O.N]Ek�PG�m��|���t4l;7��ݗ�9-�A�mF6�ݐ�˼k'�t7�aW�܈b�{��M��Ѥ9��Ne2���Ιs'K�`Z0��C�����G5����5U+u1~.������8G7�%!Դ�}�������y$z9	}��k���r�«����?˼2�����!K��U�(1U���B@%i��̍��g���U8,