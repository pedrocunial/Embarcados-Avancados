��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cЌE���MBvqN�-�	5�l��;ZŎ��lt�|���Aj�gʚ����*B&DQ,4��̣Pǐ�����οep��}^=Oq|h[wZ�"�\��<��K�L�۬<�B����S�z�Q��"QWtY�zBk�:�rK�z���i�,���SA1+.�c;�څ���������<�H�`�E��A���/ش0>��g����D�N���ߵ7 ;��),�q�f��e��/�
�t�KS�9�PYok�9����#A�,���=��@7=�m�[I�*؊s�"uA1�������G�p���m��5��{���d�b4�]��$�GՋ���2xV����S"�bnx�����Y03ȣ�C7O����rJ����d�OY\s�@U��"��]Z��ޏXI�/ V,SHP�P�YQ�wWS\[�($�n2]��w5x��ޕ��N�v^w8��w���D�m�!�#z�[
2@1��Û�o��}S2��tF���M),PQ;�=��?��1�x澜g��wWR!�u,�=�L��hZ2%��w��(�޲E��h�"�4�	c��yq0���rִl���VQ,s������4�г��^�,`dn o��2#�1A(�S�O�u�_���6��7�BtS ���9���aKoWv�v�+�M*�Si�_ꮩ�^C�́�Q���7�I�2Î��	�ޕ�����TOn�m2m���# �85����X��-��f0i����Җ����3a�v���%����X|�d�h$������Z:�L�)����������m��}�S���㣞��-̙��̛��3�2΄�$�@�["/��+��~m��wO�u�E?�j3�"�¸�G�ƣɺ�T]F��	ٌ���`�Rӥ.��G��N��w�DYI~�8IHǃ?o�d�}��H�/�$����<�3A��6��S	փ�憗�J��5`
!H��wb8RO��o��X�!��e�&R��.���1L�V�.Ry���8T��VD�����S�H%��
Ć�_�����ae")���
���㑺�cA-�>Tp���k��CX$BQ��,44��� KF ��6��:3��iwUq����_��"�[��Ђo� YrOo� �iS'���d&��i��)�H# 3 �u؍��ƒB)��s]��<������Ec���a�
�Y�->�Q;�x_����~w�'�7�glג�*���À���a�PB�Vt�UAt������%��3З6:�D�t���l�$N&Dq!-��26ֽ�������LF��nj{:�L2��!ko���k�5����_�n	���J=a���zQIb�o���F*����7p���KV`qm��(�Y��NR*e���F��d",�v|* A��$<A���n���[�Ì��r��]c09[\~솕���LP
2+M�"�9�XM�M�J��}2U/B�D^~�ӄ��(ӈ�5['�
����#�Q^�6��.왞���{�0ĪT��t�c��ߖ�n�-k��}�I�
��rʄ������X�SD�:	e�[ˈ��1ECs�ݳ�r���tM^=�)�%M��c�@�m
�MAq�=�ز�&��ٰ'�(n�:�DoE">�)�W���.�������i�^NVhĢy�g���v%�k��
�ˎ��Cc�y���)j�k#w!��t�1Ie�=
��� ��T��>��q���eH��3+��JP(�7�F�.��t~|Y����~�q�%���.K}���W�'9��7cYΆxz@||<�ׄ�ɝ�ͭ�q�1*�D�㼶�f�1p��m3�s���.0ˡ�bc�H^��SDO���kx;dx4E����s"�9��G=AgBm�wQ�F�F߿a�O5�[�Go]���eu�|�S-p�]j&����{���z��������)U��Z�ۄ�v����Jxf�>��]�W��P�q�)��R�NqV5�����LFM����g�H&~5�(N|W���,��#���ZbP����g�Dxy�.:�(�a��]�R�d�\k�t��L�1Xo��.U8��K��(�wݰ�P�8v�N��I������G�`�ܹS������yn��É[Y���X�SE%f�:���E�Y�.+�� �1�����݆��rzΡ[�p���ь�v�(��~	��+°��1,���*��y�N� ����),�s�CO'PSD�%���c�����^�.�v\���Y�("?�c�/�뤃�
4d//6��P/��jx$�H�g!�F}͂������_�o�xп�׼h�������R�����(��xIZ8�B��a�a0�^�y<C8��I8�e��'��"�sa߱M�ƣ|�+��YԒ�"QN`�}��Gq5RqFN/��N�-nz��a��OK����]��H�qL�ng?�v��k�W�ܖꩊ9��3<p�Uw����8��(��y�wC�H/(XE|�5_�6k��>$z��B3���}��Js�-����I�ZG���N4O��i���Ckoh��s���T��I,� �������A!��ڰ�* �Y���O�g'������ۣ�;�R�=�y�S�����ݿO��`�vɋ�G��.��\���Z�d���@ۼ�Ŵ��X��������7�^¤�;�j�Z5����c�M��W��_������=?�u+	���{8�����[� ��C;���,k��ֹ�(F�ǝN۶�HՉ�r�R�LǶ�M����KQo�~֟�ʙ% �O�bM%���_
�2����r��U��m��V�Xyu
�iqk��k|���\e��Pq�mq%�f�5������po���˻'������2�d��/��JsC�Mjf6�ul{s���p�AᵼH�s��h}�i�Z��koZl�����������d�`�˳4��n_mL��`z