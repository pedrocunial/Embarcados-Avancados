��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cЌE���M�S�tw��e5��q�QA��*�t��nC쉵6u�Υ�p���B�*T�Ȩ]��}�>c�;b������P|�x���f���	�����ϰ�!S�5�"*5k�qB�}^��׽��G"1�}V53�smmу�5�+V۽ /�в=�/:�l���6�4�,/�-n�G��mǷ�ʾ8�{q���}�h�,���,�W?� �#(4�m�S_�|��f�Jx��Ai8���-��X&�<���8����+����`T�wjZ�ϒ�p�.��޲lO@�y��:��`W0���Y��ǽ�ݗ��I枍f U�0d�v� �|�Z�� lϘ���pW�� %����md�ł��yo�y^����9����>I?��ŊD^�@���n����C
��Et������	���Y����׬�^�ǟ���*���
��ȭ��|�ZF{l��a��Ə�҇F_��Ę�|EO��X@�S�Y�8�klՑ=HR|W���Үr: ���/t��{/*�o���Y�rI�f*E�o�s~�/������<��*���:�MQZ���/<{.�d���#Bf�&�4`������n����:� (��)y�4� ��{��ʳ�k���|��ru�0.t�WP@V��n��Ռ�#.��X���0,j��Y��!��vQJ�/n����� uFV�w���Y`)��>�&$E�K��ƔuQ_�TGL��n]^��� ��W���Va�_=�p�b4���uMt��������J��bY	�e.L��/����!7�C��c���ռ��&߰tD:t�v�[Y��灴Z#��&R˽��Z��Q=�8Q���%p�҂��
<�&�p���lV#�x��qA��_�oF�Aw�����*򦥆�`̧�|���U)�Z��j5!O�}[��K�o�S�� ����Ѣy?$��r���QnH�eI	�w;��q��=����(ǺC�gڭmY�����>'8,|�Is�1�.u��;'�߬�m���M�<��k^]���D Qܤ���J0Z��J�Q�Llx�_����;9f'a�p��r��f�zF2�ӄ7)��p2��s#��j��oY� Z�hm��/+���!�ne��J����^�1ي����(�	�O��iMr��/~Gu��!�Pm7 ���ꀤn��'�j/w�}��-����Y�9�Eg�}����u?ҷ�� $N�h&aB�8ox��M0mu��w�O{�Y#��i�������54�[�|G�a*�IM�g�����I6��"�g_�>E�n��tRi�Zz��"2���B��z�_��:�Ѫ�%g��V.��QH|0�va�߀�n_�!G�pTT����8.��W�1��b��{+E�
^�}�$YK��0�SI_�w������!���l5b�F��.�t�-^�?,k�[4�t�I��m�7��q/b]A�2	R!1��\�>{t��j�йx�e���3��B�Pݩ��OI�O�����W�^q���Eo���j[�6������,�Ya/irT}�0Q�"i��za䣗��(g�_�=:$�]�B�]Kj��x�\~�����yU1̹8������x҈8���kU��a��g���X�/�*��v/�3Y��4uCmE����O��m�N�r`�zp�1=��ur]�����-,�'pQ%�r.�	���w���G<�+��LQ�R�=o�r0k��P�����G\��E_V؝������!+Dmꬱ}��STb���1��\����*�ɒ}��S6zs�Y[�W��f�pz��{rK�3�
�O@<���E'���6��ģ���p����n����PC�6�x�>$a}���s�� (�q?'��Q���u�yx�Y�OF�������g�:�28=@A��U�5�7=��)W:�+'�4'k�f�A��A�{��?N�Us�Tv�[B#��-��^���v|=�� 4�Hi�d�p��T)?.O��\W`������k���A�lF�kR�6H�k�<�ҽ���&��ׅ#ʺX&��A!z���u�Dʹ{��:p̉�ް�I}w;HAg��g�I��۱������6V(������S��$��{w�+�v��f�x�v�eW%�7]C��8�ܶ'.�JR}ii��Љ�|[DV��e��w>U{{�n��\6%Nb����:؏h

�ǸP�{��>��D:����3�9�r�c ���eu�%��|׈�����:��%H$ez�UG^�8�������ĵ�C�ʷ%_:�+�� ���o�\$ah�x?�+)��5W2�V�@,/-������\�Bl�Ԃh;�H���e>LC�T2����ų ^�Ͽv:�;$���!Zi��mG**H�n�
0�\q4�>&��Ծ��t��IL����r�v	�M��D����\�F�D���uh�{l��~8JƗ�ϳ�A�!|�/�Q�Ca�<D�e=ys�xx�6����<���B��Z@ݯ'BJ��<%�O��w~�FԦ\��E�1��c�B`���i�)SoU�U���*vZp��P��]��do��;"@-"A=�I8��5�,�$i:�fj~ۆ5��P�Z��UQ���׮-N��V��rL�|��	�lF���Y�G ���}��M��dl�3����<>���+��h���h��Mk#H20�p�t_Ъ��K�h�����Á��J�TAck%�,7g0m�s��l[�*?��<��i��M�6ަ�6݆�ԧ�w��M�:��BʜbO�c�^&>�sM������<����$��������׼Y�I�(�jiD�s�ً*���25�<�ats}�5C���)&
��p&�V<gV��h#���K�kb��X�uT^`�P��웃s��T`���Pgg��2Hr�-�V��jf�4i&r��qqZ7����3��#��p�9fYhFǗ�QDT���ds��Q5����:D	��׌���,�� �Q��6v����O����lY�C-&!򿷺�ђ��#�	
���1��F0�ڼ�~�3Iy�
��i�z+��MO�rS�ܺ���O��*�id�yI��K=�*�̝�V�}�=�>���'��ON�s.�.��JL�t6�E�TX�Y�P��Xޫ�-��{�� 9ݵ�Y���EE4�/��d};��n\��r�!�k�n���R_����1s��(;E�ݵ+�+�\󂦞�.���h*a�����c����W�+�sRH~{�T�y�ND��n=!F��Y�ɾ2$PẾL�I�����/�>B���H�8V��r0z���{u�Z9�����������P�S��S���C�"I"�*��?�O�z��
�To�pi�ZE�C-C�~_�T37��;�έ�|��b��^G��Z�?p��Lh+u]�`j�F�!RGhl�`����ܭ�*.2�m�f˽����rj��-hCP遄�9/���D��>����˺n��Yҵ��Sq�����)Y�tx��
4����Vh�hV��~"yb�qw�a��&�d����3��KF�z�m���:�6|$����jn��T�o�Ě*�ϩ(l'S>��V�H�č����?��!h�M
	�]鐶co�Q
��)��m�b�ONʗ�%	@�X�m����=�Q���~��6LcV�z��ي)6ɓ8��?���i�������e%VI!t�4knEK�t��n5�	q>8��P5��6��!r�AkDs�8��g,�<m�cժ���~�߮=3���2���r"�Vg�j�y�^|$i�/d�Hb�k�L�eC��O���L�fS�<?�P���R�x,_~����w?��v���Q�.Q�!�S�Me��㼺���S����r^��ӅG�ʧ>h5(�Cy�Bdy��rDa�:�g�ZXi�ز�>upd���t���.���N�:k��'dQ�!d��;�i�0\�t`Hvy`��+<�k`���XF'�-��z�yPH)g%T3f	v3n�}J�k4~��[,B�Qv���S= ��G��|�1˭��
s0Vq>��:�P�+�+r;֋�*���a8L� }�r�(7+��I��Y�aħ���ف��w����.�O �v����[HW8�/O�]<�B��_D�ůR���r��$��t~Ƙ��hJEhO�ɻ$�yK�ܩ&4��&�����Y��g�3i��^������LV�C�;|��8�k���Rg4~���[� j'w��$�y���Lo��\�-ѢɆ�8������W�F�!�(��q��l� �,n�捼�BW�� �iYJw4���Od�e'C6�"c6PL�(�8Zi��]� D�N�g���X\�"�!��b�]Q4ۜy<7��%^Gt��]��)E����%�x�{��T�N\��X�{a+8�Ww�ȏ��y�4ʬd$�p����/�K�ym��DuY�B����d��m-0 ��3Q��V�͕�"�H��`��^m���6SBOn38�Kp�\�4ius3�ot=/�1Ʀ�O�8� �����bmz���G}	�Cd��� �<��ܮ��}��T��l�{
����`ٺ��H�:���T�5vɶ�@����0(�i���J����Ƙ� 2��v{[q{9o؃m��#�Y�n�������/�+��/
$O����3yd_Y�7h*so�{��=�6d��'��hr2$s��N���UT�P�E��Q���Gd�<������}� ɓ�F����]��{Ǟ��	a��`���r��N�E`�FBZ6�ޭ�{hw�����Wϸ��±��~	 ��xf.�#�K�QL�*�oz�ΐ�r���AQ
|x�OM5̌%�&S:�WSv'�'	ڄ����~Ѷ���(X&���v�\���r0�Tj=�����]����c)�M���9`\�6�gN閑�Y�3��V��ND�6�5x�˸[�R���<0V\�9�.��a�]�{b�f2!s7B��e+�O�(�~�Pu�G g��v������k(f<U��	��z���<oW e>I�W Dw!�HbG�/���eVCݑ�5��Y�s�:����l'�I}�����e.䔊ƪ���+�j�Ẃ�F���?Jy��i0i���h�*�E���|c��4�_4����$?�͔�WƂڥ"�f�'������3u��cQMo�'PH�Cp_���2�H��)���# f�A��S���]vǲdV�0���4��C�Y�(���L�)-1��|-PO��U�����s�[�����]�qG�e��ꅇ��+�WX�*�L�`��"�u�-�+3NJ�a�ޘ�dc�Q���݇�ӗ{�
�X��y�L�/K�5��tH@K�3[��fi�����Rc�\��1Ж{R�~���]/h�Aϭ�ᦨ��\�q����S���x\�+6�����S�M�/;c�Cb�a���ۃ�҆���{�f�h�������R�'��~�^�.!�h�f�Q�� I߻�÷4�j�uJD���o������U�jL�5o���dx��{�-/��Fn&w[K�F�h�'���Xu��6��5��=�l"��Tc��5�-^��訿e��[~�$X}���'����$�i|�oa�T�@ܟ2 ~6��ޫ"KB^�F���h�o|��[0?����L:-5HsΌm��ǀ��O���z���3�WOoNs��b���L�L�v}t:0���ޏNZ�����t���s���n\�n�θ"5i;=p"��ǬzϺML�8\S�\��H��*�_�~���)�7@�������`ݔ
&�)(�@f�4Q�+�;ޖp�T���Iӓʦ��u���#Mr1ՠ�Ti	�6��y���4�EP��`����1k��qw�W ���X��l��1���Hh�8�����-m3�C�/Lw�H9Q,�����-Lݬ��9�^atfoO��,Y��y��pU��	}���`,�j�쬮�)�,
90 -x�K��+Y9�3e1N0S�Z�rH�k�Â��ilӜcj�y�Rɫ�a�Q�0�XQe�d�����A:��r��LzmGD��k�+Kk?�,g�vu:o�]�՜�L���dّ��3��y:ڻ���؜�����	k��b��BB�E�����������w��w��6O#�5��3i��G�^h�|�F"��J�����*~�|eN;�{Ը��Y�g�ΙҔ�f�/ �c&�6I
�E	녲5\[���!U�:����k�ү��b��st_B��k��`Ѿ�k�b�.B���2��
,�Ѝ��]AU઒#r�p1֚��,�m���]��?���:��Mr,�/g��1`[�8�̧_�h%O�;��[�/y$l�t��^�!x���0�-��7� �N]GJ��M`M�Z~�9�(�
��^�����q�;mY|��d������r���/+��m?�;�;�o��}9��;���b��g�{�K�-)=ٔd���Q�l�w�/����<oQ7�g�����?>W�B���!w�I]z�e/��q�����5"����'����j�0��I�C�i毠`�:]X���<.�%W#�yr�}'?�ck%�-=��.�MM�dž)p5��r��`�5-���fdD}�U�w(��֯r��o�H,%t	�÷_9�	�#��I��(&\gtL�z�[���Ky��ɥ�Qc@�i�C�1�U����)���)3�Mx� �+)�<9"�����#5�M�M�Mf�ҟ�/h6P)O�/)�s��ywb72v��=q�C�xߴG�D�#6X.�Ƌ�)MJ���,T9��=�s��H���")؈WP�;Bϊ��f=ץ(������$��G�\}��	�~7@�<��s6��bh�|͇�CJ��Ѵ��zA�a��_V���jwn����S����OB%�V��jQ�;��M��m�Y�̜Z)��M����K�|/M}G�{x(�O�I,�A(�i�]�K&�U��V^+�����Ƭ������ᄱ��?#��n��T�gy-�GHFz�s ֶ#�/Il��	N[�X�Oe	���or�v0Ë#OR����+���$ڹx��x]����0΃��>���GD�XY��n�Z[ ��6�Ĭ�g�
��of�<|� v��Tyf		Ǣf���t��D�~?�&M�7.NS�����]��ʫyX.��
oL4�+�kW�GCI\��w�GMo=NMi_��͘q��2w��9�k�p����/d�f��Pw�*A��7х~���>ڲ|x���@��krX�ƕ�/�� �R,,z�����)Vׇr��V*ZA�x�uQZ��\�2dp��Ռ�{���*�ꖡ�򟍪�W�=h�Cr��Z1��	�B}�\�X��'X> �߅�� ��d�Mq��vK�{t=��*�U!��d�r�v�|�� ����L8e�c���<4�Ԧ� W�C��c��-�N���g��	��-q���G	V�{{�����(T���t(x��DR��:Y�x�J'�T���#q�/+��Hi���oO�S�%�*D��%�@�@�m�񙇍�M���?�Z�.��L<�Z_W�f5�ޕ�W`g��jS[��)@���"�K$�<ܟbz�m�����{�.ƒ�<y�A3��+<���t�$����b6��Դ����T]E�9\H�V�rp.���b>�GQK�4Eȳ�����/����.����՗Kc�������<�)�_M�Z�(�s�)f?h� 鹸!�5�Ӿ�̡��!��� .�q!�~�7$F��;bg5��x���@��4�U"�>�ʴD:��:!��B��0�/�����q�K�vX�Οs ]sR��\�,K@��.��N�r������[�֫+Hv��i=��q:{e1<���tl.A�C;@����П%]� 9��X��Ν�e��\�"�65��H_�͵��n�(�|r�a� �Ϧ�6��\jm���?�����gD���O��:P8�/$�	���[<qX�SP������������@������f�)�I�I�p���aDF>���K������Ӂ�vŐ_�X�����Ш2ïsJ�8����Կ�*b�E�̓[w��D�d󰝶r)z��k�o�S����^���ưS���O̊��3�b���>�@KRqᷴ�w�Z���9Iy���k�]qS"�Zop���ə��ԑ���X��=��D�e �:D�ape�G���g~I�'�pR��/i��l�x�\ĮtU�갓���0�.	�7Eα�oi`������r�9���I+7��A"�Cz����>�Wn6�p��(�
�p��� t##��.VhP�;�/�1�3.��7��+�*S�M�R6r��<U�h�,�%��߅|o��H�PZ-YJA����:1y�Q�K�����8Uz"�j�;/a3�)8&s�m�i��1�.���������yb��]!��]��\�Ij�83�D3�2x��TLxv/߄��|g���0(�Z�@���pD��^Ρ��;oD`;���hzڐ�݊_�i���(%��;g|[�_���ͯme;[�c�R�:/_]��r��&�Ԡ��ꀃ3�SĶ�Y�)���H�����⏧����Dz	v'b�^�s8��#�p�Z����~ܭ��j��H�q�d]R\��3"�E��}3Kt�L3?�o]+(�w�N�i��^5�c��� 4j)�2%]\�k���w����T��+�����OM����ך�1���c
V�n=���~�I\�g�?�D�} @5��?��9��?���C�
(l��&?:�ʭN�XD�?�GJ��bqm�x��#j��ѡ1b�j�%��d�tR����.4�w���S��m�����6 e�!����q���?An ��D�'�Tb>���%u�.�:0t����� ���M��?B	P>�����!x8-:R6$Ցsyg��t����y�0/ʞ@���>�����h��6�c�c��ty[�7d;e���xy�#H�^�7���Xv���%�ԣ3��#P���,�0�f�
��fm��5��c�j�������*C�"
=���T�c���0`|�xԒj���DS�R�R��S2y�)��E:U�w�"$dd{�,�o���k)����k��f���Q���7��gD��O�]Aj8:���g�?���tG7s�����`	�35&~���k�޼f�2�U�O�����]��ln_s��Y_�M?L�4Z�����F��t�h����@$���7Wͺ�����_|�L�A���=
{sh7�~�!��pr�Z�@Vl���KJ���j�J����_���{u�����q7]����d�F	����b�&?�t�j���o�|�p|�����̚K�G"Į�|;+dƀ�� u���C<�Z�	B�I�pYiviɮ߈1|���n{tS��+�_;��{�w��)v���%�p���8���w��u�c�*����n�и\c��M������8ɴ��)�s�n�
"a�U�溦�%d��J����}�5�?X�B�L�*.�ܽز��U����VfK�a%%^d"W�Zɾ(¾�c�<�ő`�8�މ�����H��D�d>�J�w��I ��t�ЈhH��L*�y��"~NvP��+x�T�D��8�?��)r����i���#���1��c�I8������i�<�90��~�e
�tЄ�Yc�ï��=��*�W�>�N�]��8��!{�M��"����� $�Е\�l�=���V�=ZBf��'(Ҧ��aۘ���|D/,�/�
ox��քߏ�O-VN�h��F�� 06�"�i����&H�TW���[Ԁ���<V����OU�F�Dۂ�-/L�{.�ҹ��,>+{(��%Zs�.+����QT˓Y���ű9���N=�)��洰��`�� �+�`,�!���-#	fy�+fpZj�W=���A��:����`��@4C�Ex�h�'�����~�[��O�B���vr��o1��3��)E��R��jk轳0Ŝdˑ�l�Z�i\�/r�P|�M��[�(�*k)��D��ډ��뤷���yʧ��=���Z	¤&���P׵R����:.�i/�0���-�������y�G`h���耀�ckը�3�#�g!.

��W2,��Ƀ"r�_H���J����:'�O����9<�L�O	��CC��8M+�/6�k�Ǆ* ۹	A���}	<#=ɗӈ� �Ld�Q׮����F���|��(+�<^�3WI����` ���~�N��b���kK������lIxX��	���/
/��r�S�7!�k�fý2�A����׻Z	)��-ֽn�sB�l��z����9ؔSX/QB	�zUڶ��?49"��\?��b`���Gj��������&i���- �D�G.�To���j�����t��h�.S�cA�^��NuQ�K��%3#�����j������a3�u"�*�X�d�SJ�藋�+�D1k�>b�c��ޗ�ǃ�cmS%���_oPՓv��)���6��ͩ�M� (�r�Ȋ�T�wds�>^�
YՙAK%T[�Bq�M����7�N��g�����k�]ګ��8͐rP)�G�e?"�h[THQ����e����m���P���7]�H5�Yܒ=��.�QH�7I�b�ZZ9��r�+z"�-̑�� }6�Z8֔0Q��lj���M���pY��s���*OPƍ�䵶��<&�tR�c�-`��j�qO�C���Y��Is�(�*#�¥� @S�X7�=������'-4
���LjR��nv7�
x��Yɬ�1��T������U���;X�:sLBL ��݌18o	n��=��׋;3V�Ix�K�d�]�����g�q��(m$�\�A>�@b�J���i�ْ�o|j�*�Ѧ�2�9�.m8��j�Ft�sW`��$~� ���~�Xi~�M�k&A�<8#O�jv��+ʠ���~���b3��zc�	�1$�I�y,7����~��r��v0���*��; MV��~�����d"���c����iX	��AXR�t����46���SЌ�יg�o�Ϙ���zv�Qn�%�T����s�o�u��)���N��������k!��\�I�H�RoʠШ�h�ь�*����Y�̧)�[�~g>��F�l�����o����ϓԎK�����E@A��'p'c��<����3�8���������^���ǩ�A{�����e��M�����Nmj_Y�sԪǔD��Jc����_�t�\���T��~����X��ׯ!��V�PL���;�O����s�'�&G�r���|>�f��y��]9m�^
`� �� ���@/�њܚNU�c1+i�ދȺk��q���J,U��L�)*� ߃T�W^l�(���Qߛ��7�9r >n��y����%;��	�y���(䀕$�� ڸζ�Eִ�e������;yehCI���FX��Ռ�Ea${����ǌ�r�\4%�]�4�X�*u6�mNA��ګ|ly	���&^,�h�Ze�$[����z���S��%���]��b����nZwQt��;����2��fm��o��ca/G� _	�� �ݶ��R��.ŵ�h���4,�m/�n lБ�i&����j�;��Lu�SUݏ���c�s�^RO�Y��:<Z�����+����y�8�d7��6��Ѽ������"��> [��_-6���
��Yp�y�*���$,��)RO1���Mq�����034
� �:<�Ԍ#(G��'~~�$��97����?���G�d/�!�����Ǒ���?ߏ��^̇M��ADś�����O��3���}��<�i!�p0�FS���3��WQ��g��?+�X~�O���|i��.I,։�/�0?6���J6C��(���έ�f��02�1M�e�4����� p�����uM�	�];\��/��?�w�Y����=�/.	�N*ڼ(��D��y�vD"�Bt�yÑZ����;v����`��O��
\����z����w'��6].�����LͬA/5#�ɕbC�t���`і��'�Ǒ渧��t���?'��FM����z�e�f�V�e ~�[��N�-F-�o��b�6҇h��i�7w��%Y��'���T�X�]��\ns��̹�W��"�;y��`�y�U��SU�j;�1����?�X�T��탶4 �<��$1P��槮����r#��|�����0�>J�9W�
{b}�7V�!o�YzN���J!՛�ۯpI�������9w�?l�vb@.C7��*'*n(~�Y3ۃ��>��T#���D�q�s���ȮȔ���k�u���^�%������ӇZ8�x�D���*A�_�_�T�*��f���m�1������~NZ�O5§e,Km�S���
k_�d0=�B� M#-��O��D������	����ը���⎦���W�����\C�Z��LK�4K�o�?3�)R��E@��iY�w;c$9ޝ��w��Gs|�7��s�$V�Y6Wu6jkڔ��)����H����<-#�G�!^CD����1J;۶����x�<�?!B�>9�(�d�#we��4�u��0���3�3`X���s�&��Jv��ڹ?�9x��<�d/8ޏ+q�$�n�ϊ��|�/��(�Kd���-B��O2��!�yT�����m��YYlz"�Ϳ���y��[M5G�U:���-�Z�Z���� ��A���=ػE����(%Khw�+ؔ@	�C�����[Y"���d�B��Y;���& ?�ɁI��Y7S�%%�o�:1��c����$r
V���r����o/+n�iҾ���`�R�àe�X{*����^�i\��r^=P�Ԫ�Y���_J���@���~�f�V��U��W�n�C0)~�	�	 !O�xY����N�~%%�����ʙ~|���o��WKx�䣌y
�RV�xN�}^�nŢ�OڀDJ�'�v�H�ʈ_Z"d�F��-��Co����Ƚӑ��N��3�?�eU,��׵~ԁ�����3I,;^��J�������r O�=�����?J�SS���h���F��`��s۩~ԓN���[KW*&l�C�O,f��ViG�d[��x�R�co:PR>��䕟RL�����	�IqB�g"���UL��(��2(�X��6n��:ֿ�>p�Y��^��a�JC��r]:D���-kʑ��+_Bl'y:�7(�~�Nz���
#¨w]ζg��#�zʦV�9��<д圭�Op�lQ
8)�@��@thL�k
R�Bt7پ��_26R���$A��Ӟw����>��)�%����Yg�;Y�[��t������<��A.��k�$�#��Fi�|��(��B@e������]���Su�~#ì�;*@�,Ո@F�u�͆SmL�����辆TA:�A���7��]���َ�M�\%��_���Z���* W��I�׾�$�H/�pSա�ʈP@q�8�z;iM:��ᛢ���̢�ר
8 �pғJ�9O�t�C����?��$��ce����xo��ݘuS���f@ (�G�э��ҫ `8�mY3δ.���]��WFj����e���g
���h��2��f�|�����{��>x-B̽,���l���,)Q�>���ԥj��&�lvE�H��7 ��<�l��	��[���#�ȉ�0�^����$)����=�Ge�c�7Kƍym����5��u�)�����|��7�K�<)}������A�y,'O�A5�p���H8�"��ٷ�檼Yz���ʌ����_�KO�̛�c�U��^V�_;Ɇ>��j{��i�t[��2�e����2�z*�K5��QS(X��C���� f:b���mE����2�_���*�uo�r~n|��U+y�w�b�*���w�:�����_a��-��$�z�������$wUe�?�����^��)����J.S�̤ �7Y2Q3�ep��O���	}��4��[�Ff�HO�c@9�&��,���C)R���c�r��ޱ%��΍+�i���H�э=@x�G9k4����p��!X����"
���s)��z9��{��*Y(��tԽ	cth��w�g=6�������A��э����"�u��=C�
!���U��V��QA$k�o����YV������+$S ��X	{���M�z 'r����"�۫���O� �y�bH�A-�_�q��j"���p?a�%����) �,N�/��+;4wi:K?�f_���5V���N���V��[;ƽ�3`q'��F1�i;������#~-���Y��[we&"�f@�Ƽ�kCl����dw!�!��}�m���q��5v�ۍ/O�E���/�s����nσ���4ўy��οfg��}H�w�m6���(�&��^���o��7���K��g�}�n��폠�1?Q������.ev�q��P!�M��,`},)�v;C��K��	���(�TR��@�����	X���u�Rǧ�����%S���=O�
�/�Y�;E�1-��M��i�:�������Wl@q���U�o�}iO)-c�����<��e�ѩ�*]����[�aR�!���r&�]��!��I�#��Q�|.�s����������]�P�'�u���p!��.¿
W��2�a���G�K� K��..g����}�f�vŁb��f�����9RZ]wR��P����X�QT����,,��ѨZv17�K�{���ؠv\$nUc>-U{�6$�o5�1�>��Y�������+��x{�Z�������B�v�϶F��nUb5�@��ŗ� =/|�Ӯ���:d�S/��s
�������B(l���32��>%�o�ݜ��Q�� |�tU�WYm�E��rs/�,㟈�����k۪� Oy�w�����p ��|%�W����=�5���G�]	礢���S�A|����ek�\m�^"���S�d0�*Й�>_�rco�G�U�5ې�D '��aK#%j��XB����}t�ţ���yW�#�o��/:�����b�mp��P'|��H�TQ�m��3J1��|7 9f;�K�#�ew�y: �;\e����SE�������w�w󨏌tɧs;���Nޱ�0E���+���rYEr3G���[��m�I9�����3,���Ce�!s�XE�)ғ�3T�b�=9�*h�s�=���ԫ�fu�]�g��F�B�֋j5`!L
���L����1jH�@�g|�a@�+ !#=�=��[� BfeZ��k��Jé��G�C�����g@�w�WGR47��A-�c�JJ��)�	D�3��PQN0;��Y�}}��졷&%&.���0�;Y�LH~�˺H��_ �6�	� )u�3yc�����Y�����V��{L��'�M(z�3���=Ty��àd<�՘����+��P`J��F�DI]���'k�Z��P�UӋ����7�^�N@o�ƖOu��jX�)�����R{M�kr2��w�
�=Aq��ZZ��H\�(n��Yx����W��h��D
}s�@_/�QztlP���?�u�ѣ��d�ɓޛ�ݿ��ŵ����b>|�j_�mC_���Yh����q.��/���}W&Z'�gK6��!9��x�'��51@�of��V@�������
�-3mB���lT�Vj���w��3���/[�5p��{���/�Ҫ4r���D��VE��#W2�.0Ȋ�u�Ġ�������d��w��v.:��8n6$<!=a��f���{�(��[��ˎ�LCK�o*ۍ,���v�[�T�b�AF�M髹��]̧1�$���j:�ą�d�f��o�`�ޢk&g�&�"5uF|����W�p��Z�2��}�k\�:���lͼ9�1��S��H*���c1n���/���T��G�iAZ��kp9V��� �v_PaՓ�S���� æ������3�^W�Q��!"��Z���/͝n��WklUj55y����e�����Dҗ �?}�F-�� G�\3���m���e ���}'���7ƅ�~3��w��v,x�� V^:O�=R������~[��~���������.P_�"{���*+q��xp }���L�_�Cb�,/y@��ő��l���?|���\Dmv;����ʃ��Z��7DW~ۯ�D�FT�K+5�(��%qߒG
���|ٯ��LWO(���d�j��n�l9��Z�*���,�%Q=�������y	�jo#�FR�ri���k�#A��$Ơ��km{�^f�i��+1@�L`�g�vK�my���'0m�o��D�Զ���6E?0��aQφ��8�$wA�(B�K��%]�]ΚO��`I�&����<k��9��@I�Jۃug��\ӳD��ILA��(x�PLc&p�ئ r%�$�Rs\���1�2g��΃@D5=��$�WTd#l��'�}�A������P3pMp��|�&�[�,�����τ�e�t��Dz�\�W��є���߷��Ӯu
����`�?P��� 2*�(t��+r��Hr*Al�%�x�NsO�)R8d0�i�Ϛ�I�u�>=1�(r�৒�vPI��#��dO����s�OŒ�^��­0^1��Pb1+�mGmV���|3��2�`8YH�}甎��Vt�<n$�ي��hh{l�Lk5�����&��H�W����&1,�bj��9�����v�IB;�$Y�*ž _���_t1������و�Hdr�w��F{�;���l&���?���MQ6C%��;	n��"q�w��)��-���U-0��S����R�j(@FF��HE�>�L:-ƥ���B���Ձ�c����;y��
q�V�`#wkF����~u`�9LY@v�	P�hCjxejLÙj�e8[QS"t6�G�`Y��FL^�����b��3�m �I]ӟ���4��8�!�i�D�_?H��R�1�J�Um�cg{-xY��}�V��BU)�gӉ0F`2T�&�7��KQ���R��߼g�x[w(��M���J�����c(��fґ�@�! T�����3�%Op-:+���'�$1�1s~Y���/�C��+m^�¼PB��oE)�xu��G��N \ia�Ъ�h���ՉU�B��v�}�2�"o���R6q�Ez�������e�d�