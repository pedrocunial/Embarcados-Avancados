��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[c�Zz����!U�=N;�$5��r"��bxl-�w%6�ܒ͆,��=�I���$��ۍ�+�$����y��h̴���� c��_2F]��W�BZ��Ȋ�c"�@J�ԳXɡ�ĽM�=�5x,
���H�uh��=����ܕչ���%�:Q�5l^�)��l�\x�K���7\Һ:S��M؍d��9
v6r�I�c�n��)ʹ���>��TEiD� t�
�������P&+�'/}L��4(��ż��v��3�J��2�7#�~��茱j`�P)U:ܞM�#ni!cW^�I�$U]���R\%�iڜ�YUJ��~�A�x�N?�j��_��S��\���{���PJ�7���K{�A�:�fE��F���]���&�Э�T��zB?y�p��Y��<�h��>ְ琡U�F�֌����'�UV�wٮ�|�&�ޫ�\܎�f�UN� ՝D�5X�b��X�Sɛ�s����<!��@�Y�oam��,v����1>2�Ѝd���=��m��Qy�RY�`�d�#y�\�<%�B��A��oh�����-D������\(|� �&Ѧ��t����/ |�W|?���Y��w��(k~�t���&(���Bwbex��u3o�柰'��u��a%��`
Q�ݧR-�҄�� "K�3`̮
�h^��J�����4Vc��`��N5Q�k-�;c��*NoTS�Y��O��ubb�q�N�a��*� ۦ}�����%n���q+�yQ�bL{����q)����%��RX<ǡ��W�I�Ʌ6y���U�Γ���S�C%�J���!�(u��;߹�p�}��Sӧ]# s�}�}��nb:���a_�%4��<LF|��Y(iT�i��y��m���g�s�b�p��+|�u���u���Îv],�d
�I��[�6Ji�� D��6��-ڼ�|���5�jt���lC�c �]�3�ѳDS@�F�B�eGP�K'a�U�j݌_	�d~㜤��eA��J��H�o[���@��~�Q?;�%��'�3�P#'�C��؛#����'�M��w'�������5�g���d�#�d�A��竅�>�#��]��Y���i�↖KR�9ֿ�P���C�fRS�\0]�-�/U�Iwyj���`�iw}s��h��'{N�yM���	�d�$�����x��������ӆ<)�������衴�Ta�QQܢ˃�j�ۏ�i����r��@��y�����^|��^�n2Y8���H_���˵��ZDĮ����{�X���&�OR�$�W����f�nB�r�C�qTe���yj�1c�L57�.O8��U̎r�0*�ƉM<��%-�J�m��E(\��д�]��G_RwƆ/H#�!�$��S��!{]&��i��:��Q�?q���8΃T�y|�hxp���������ߝD�QcIL��λt�ιuX*\���	+�a������[a������gD�.H�n��	hG��I��t9��B"���˜ݟ]�UsX�}�^��]sMrR�9낾q��v�)
��]kT�!V��[�p���F	Z�cWM��5̾K�BMm*����e��m�=����T�:)�\gm�w���r�*��Vs���	�?��{��A�	���
���?�V��`��I�u?���-�{�d:�z�W�a�f�~i�[�H�*��X���Ki��� 
5�'֫x�Њ?���~���H��4�$� h��C�I&�a �
<Z������A/���Qa��0?Դ�h��������5ɮK�|��b�5Q��R�'�w��2 �}�s�0y�M[H�0H�a�,�4��qIx��mDì.3w��\��f}��Q��~6}��u��#jyG}�[�~��	GI�r��+��д*�mjԁ<�{bA2����}���Ͷ����ü�_d#Ŏ<.+-��_6��qD�޺�Q��W�W��ju���o:�入�m���`k�j|I�&=,�&w5wF����]C��6ĕ�3�C����Z��ѓ���7�1�%����I�g�>Bi�C�73&<�]k�mW ����U霟���^�%����%��{s%���M�֋Mȥ�8�������lf2�o��$+�.��DL­	ԏ7M�ve�H����;
� uN�d�'�z�T�һ�B��=H�f�'₿}lmG�6���ҚM����)\Fd�3���`��6k!�b�BC��4�ƺ2l"�e��]���P�h�73G��UC9�C��i��_5�Y��y�;Q�@���Z1sp)vv�ܘ�U:L�Z���|������E`�g?��'ǁT�ҁi�F�i�XM�<,�<By��s���zi��!�Zb�֖��Ut�1����my}��K�������7��`�g���J��ϊFEY����e���3��f�(��?<�aM$D�������Ǧ1,�� �d�3�R��|��;k<�+�k���]�rJ�(�o��Bd���u�W�p.?�_#��;ަ�-�Z�K%��봿�_�9����/<NX�y�����jք\^�9�+-S�U�ML�b�	�
I�����QUր-B���U0��i�򂮯��z�C�p^Zq�<E�����(����H��)��:���N;\��H;%�]�g����c��oڏ����������Ҭ� /��A�ѻ��r������
��U	��4\��If+��k�HH鎲��j�Fn���͍@7�?�w���V������$V'8[��l�:s����1�"2S1�RǣP�����#�T�eԂ��r������.��Z����%y&��@78�~(�so�YyE��dO�j2Cr�/`�=,Aس:���.��}�E��F�5!���_"�WgkB'>�E��R4:/Y��`�l���z��c>��}'-lB��A�#0�1P΁l�MR�L���$Ce�i��& s6��߅A�o�#���s��S�Ԍ���
u�iy�To�����2U���5��U�b@zM���2m��~��\��gW�ͫ�nR�'�)�"#�b�k4�,�zS��t�-&��:�op�}�x]���7���A���(�}Q���Tz�T�kn�+�*�E�ѱr������샿hǎ�غ�D���~����B�2#F�ëW��d���5�
N�VO��Hƥ2�<���E<Ɋ�#N�i}%��UhK�9M��@����D�=m-3���>�z�;<f��J�{֨u��bi[��w��+m)�UJ0k+S�i��H^'-������ +��LEv O�Ž���S��\"9b	�������#�� P��-=�8�
�@�����@=1�ZPFQ��.�:An�=�-j�\��w[��Z�2�E��Px����U	1-�b5݀I��&��]�R��>��m[���Dl��KS�Ȅ�o=��[���|j�x�n.���1�!��Z�C��o�M���\| r���������ͤ�+�pBFmN���3�o"��4FXc��D|��P�n�#�<̍�K�) �Ƥ壏^Sh��t�Pa��;D"��
V����Z���JG$�=��"�ry�GD�0��0���O�S����ɿYoT��P��	5��0yܹW'Z���^��v������y{�֌��B��1S=8�	m�v��Ҟ�@��ot�E��Ŵ��[���=�W���WԵ=����R��~�բ64+}����w٭�9M�4�w���~P�Z�3���b�#*�8�0V�W��V_G��N-��{m����`����)rk����ۡ��ߴ�P�O�qv�Ip��kt-��x���jH��p T+elX/���t�
�SW�	��A����_n���� �,�k�-UtA�xY�*=��zaFJ	=`�xm鄅Ϗ�L��;�ҕtL���@��#Nq�5||��q���nΙ�o�,�Vn�$,l�[��R�k�\�Y�С^�4�o�=6	�8�^%3Mp�=��H��هT�u�2':;����h�RG�e���~I��?x��#�iI�Xˤ�T��<Lh=ޣ�g�֕��@`M���0M|�+��2���
�@�mX�,D��rVl"l���j�i�B�7�U%�bီ�`8~v{���.����E�]$Vt�ɩVQ�s����t�",�I���R�^_Hɶ����ߗZ���+y�BgY�~�͇��&��M��lV�M.� ��^�����S���_UQ�>R)���CdS_%��yy]8���R�|�@��F��24Z(�0��YU�a!�^J��k�N�d:���{�:����;GE�U�H5ۻ�j��q�ZiTl	J5��oM�|P&��c�W�BC�|�8����Ơ~ T���\C����}���hAB�So>?�J*�L�g�Q>).D�_8��a��(��{��jĵ���К7�_Ґ�\%�K�Qڇa"�ۙ�����*'�\و�	]��	�? ,b��Ҹ^���A0͗y�Ԯe֌�9JnXY2��H7�o�@2�5pm4ET�V�9.�O[�C���X�e������5"��P��/}2{I��a�ثV�G��U�O|ԙ�2M؃���K_Yۂ!=�k��s��S�0�k��D�chz&� (͢�q�`w����=Pˆ�+���M6'sst���G<<����s�(�Z�ZƴBɢy뼐���x�0�Pҝ�o�70e/����B�1�������PڐlL[M)�x,.[��k���*�>���GKCo�qb�����h�S�x�\����!O�oCHv��K� !y�JUw#�L��Tr*�e/�p��aB�tU��.���X}�|�u�Mꕮ^�"��<��������m#lf����K�B��])��;���
C�����fj%i�X�@H<3�F�m}�\���?T`��;��h԰v��{�4�������Q��>�$sDD�|o6q(��gI��t9� t�F2n�'�?���m��C����Ȝ�3a�H�������(yWK���/�V��<�m�!O� Z�=4.ݫk�`�g?��}_��c/na�Pm��^2Gu���y'kPE�b��2�$C^w�/��ppX��q9��2��S��-���A{U�0 ]���)�W$S�f�[t�lX�vh5UO�g����*[��!f��"���5�̓c�Ii�n��ߐ�r�_��x�Ƿ7��T��u,��Q��d�}ݦo�)16F
IY�E���%�y����Ǌ�YR���ewb�DCWs�����9��ϩ�3��;"oq���]�M�$l�ܜ<o~�)������S��O�199�)��w���F�h�U4����َ�#p��E�.�T�ƜJ�:�4��h"����2O똴��$��妐P6�J���ifD��f�$`����wf�V�S#�EԽ�[N�1���ƻ��%���h�6lS,UeY�/BB�մ|�1�T"�{�s�~�O|2ݢ�
��4Љ|s���XDlU�@�a`����'T�Bo��O2h��M� ܣ	r�a���*��Fc��y52�?�&��v늿G8�̕ cA��g~�̵�C?�uW�g)���<v̎d�yFH�p66�睶�=ND��`���B6��/;՝��%�¢�!���c���G��-{�,NK� �5�蕃.��vR�D���@�E���kys�;�*����H���PP��Wʓx n��N\��#��
xl�xb`֯��e��o����g]e���THx+�oؽ�}&�;��4N��q����7�R���z���Ҳ�Z辯�+7:8@|�X�~�"ܭ|�n,�G:{�z��@4u�d��A^���[3Ki2ΐ��q9�}���jc�R]EƋSϤ]���^�y�uND7}i=ʶ�21פ��RW�[Q&��4
���ӛ���)�fğqG.w{u����Z�;'oq\�{s0��@qn��������H$ӕ�GX3Y PY��H��ߦ���?�+�1�H��`k�`;\]_�vG�	+����<-�ȹ