��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{hi��7	G�����|��4/���YEs��Q��H�9e���ϒ��(��t�.�?�ѩ<�Փ�<�Evj���T�����B�ݰ7� ػ�3��p�����D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[���۰/Zu�(�l�N
nk�����'��m�n�뛗�mF�觴��F���(�wNE)�U��i�ع�MyS���#7���g�/ AXW�,D8lɗ��+�")���?�F�;up�l����c�{BOzB n�1��б���ƶ�C+���_f�2�EW�"P��w@�ґ8�*;�2�p8tEt�%*7���4?�����Vo��S��޷/N=��׸s��������{���@�l��� ��ty`|�׵�xgq����#�,�H�9����H��hȻ�w�ff{�5��[(J�A@����+�k�[]") M�̡�L�q���G�#��6�5 &��9����7g�m�,��2jL~�M��@�z	"E�o��i�$C�g􋱗ի�[$L� �zj��6�JWI��``�#�5�xc�(��q~u�bl�X��c�q���h���U�&�dF�N&>��e�d����>��6c�fG\О>燺{��8g��qd
�6�KSR�c^*T��@Q{3��W��1��+�/Պ�l�CcOG%�$�$��l.�"��~-�|�  l|y��O,��zDZn�忣<�hALP*,ă5��,�77*�Gx=V��3`��$�>E(.��¿*�����>3�<C\薵{�>�V@̒��6ʆ�a��TgB/{/PpV���`�3� Cs���ѷ�~�^P5���tS�����}�<[�O{�}/y8^����Ij�R���6��zS9�ZI(b_a�D�[��ۺi�5}��R�z���$�������z܀��9;�jZ�B����ikK������Q���Z�W����@)$�UOD��w h�TcX#��АDK/=;��ӥ�G�kUL�`c��&u�x
%d����.����Y@�~�*��U�SP�U��$�Yl�"��!���v������n�s��<Ҧi-XB��b�V/���1���-as<|�d��w�m�D�L,
��S�������ŏkfB��8�֕�\�K�� Yc��a��L���)֥�P\�D�@K{f� �K۾W�6�Y��x֝O��.W�`%�.��!���	/ޑy�<�:.S��<aѸ�l�T���@�E���F�݃����U�5�ޙ�k�|)	N��� �͹����{�o/�����)T�=$�ւ�i�`�'7,�'��[��]���c@��T���l�2�R�}��vrA ����r��*��=$O�&	��}����GZ��D(���C󧭸j�g�Hel��)�H��S����#�݉�i�O�$
� �H����`�D<��o�-KDr�Ŕ���b�W��M-�&G�F@nEQ�.��*��[3�T�!�Ű����s\T���c^�d�4����$�p��_�/@��ꠔ����		��q�G�❛,�'�q�����)�J�z�F���f�c�C����&��G��j��<���-݊D��J�O��Y�K~OO�1?��Ŕ������j4�!q�w�·��$��oT��K�B�$�����$��r�~�[�4���>H��̈́�4&C�"./�=t��q��������u!CJ�61i��T[�1Wuc�ǽ g4�T!ܰDT�!H��\�i���++W��d�����yH�4��H��
�<�%��w�$�O�.v��P�&�|�9��8��]�\�|�����>-��Y��O�?�4��X����m����ĸ"�B]�I�>3�1X"�T���uq4u霚~�dU� �_N�#yկ��9?GJF	����*)��BR�Cm�v�,��lݿ���E'��t���l��\"?A�S4 �e@�!������z�;��� �0��Ch,H���"΁�>�վҮ0.�f��p���̝9!o���{w��JBa��@aB<���j�a�"C�Js�`p�0�͉.�o��d󺸝u	` ���BȎY�ȇ/�ÃWZu�|���OR���g�uѽ�d��|�1*ęjϯ,�5U-?'g��&�k��ǟw���BB�{�d-��u��6ld���a�6��L���+�x�a�X�@3��h��^�R�^�O0�/��L6��NyG��=?��s
��)Vi4�y��0h�; *��x|
�=T����L3i�����}�MP�8�S�����'�]`�g��dz���Ӛ�� ]+,�4:�nMyA-?��q��mw���U�����5Y9�np��1�t���C*-'����_U8gB��zZCS��XbxGM#���"�eG�/�>%���m�tӚ?TcR�#
�;�'L�jh����Y��� �b�kdş���r�����~n���ψ��9�v���ظ+����b�a��x�`�4o3"Bp���G��(��Q�z\���x���&��~�|܍��d��Ap��룣�%�����B�2��B�_N�'>P*	˙
�)-4ej����3]Gp�_���e�y��+�	p��D� ��<E,�&o�q%5�|K%9)���ߜ�q�k"R�It8�F�_��o��l��{�43�I�̘�f�2��3Zx��� �`��&�F4����T���?�p7���т�����
��Fӕ���2X��gF����+g]�da~�f�/���3Ӊ]<m�Ū�3*k*�A�� �|9
�o�֠���CTI�@��j��=x��u>џM���,@]��{k�����kc'�ꆠt��`�ZQ��S"V7���j��)U�.�ŋiU:[J����(\���{?ĕ����Jzb
�BB��b=ʸ�?���`��e�V�	�?�E>R����~Օ��4�	=w���fK#`�A�"ƚQ�U�OV�&a����r( 4Ax��{g� "�m�N�$�e�������/��xE�J�y%��T[m�ok��rIUM�h�j��
l�=��j�������2�gQ���'��X`��I�w� ���R���rk�%.�4(�<���R�_P�i�iǤ�����8n�J�� ��,�t��D�d�!{G�˥���-z����u�R3��iH���Oĭ%?����������%g`h�)F��*GRh����_�Ӕw�ia ����=��+�E	��z��S�8�5��+��������G1ۡ�����[�4�2_ڻ�uh�N����=�Xn98Bh���kR���{E)~J1G/i��1�t�"�>3�IUܿS��6-�*8S$/���̷ éݞ<C�L�!�cD�^Vٴw�O`W	Ч���7�n��q�\���┵rCGf"%�0Ӻy�jE��a�zK98ޠy�A�T-5�+we�W$$^�x��f��#��g�$�B��3�-�/�k��u� 0A�,%��ͼ��fL�/�������'���L@1k� ��pu]����6���΀�V[f�?F�C<�@TpVh�ne���L�vГQ�FQ�?�ּ��ѥjQ���-���'(G='wTw(A5��L�GP�/��NHf�C�"	��%W�S�P��.d8�T�&���*�Lp|��|v��M o{h+I���ILӾ�0��>\�н����(#5�;{���tq+��vvk�c�ݜ�E��R�������n�;$A�<B\R�.�ۤ$��Ԧ��.&����<��x-���3��2J2��'��s���w6%ra�2��~X� 8��FEO�C*nW��4�n��2h��{���<��Jo���Q"��(���E�Ù�<����@�����ǁ�*��T��*�������7k���`�ɘ�ά.�1�Z9� �%��g��vKee�Ņ�iͦrWmա�|HS�X��$vj�$�p���j��!N@ȭ���5%&���.�|-r���.+��zP������ӜXSc�sI�	@Q_t5�a
�|$����*�������"�h����J��p�N�y�D�V5�aM˱II����R�P����w{�cܴ�xK�e�Y��΀f�0e�?A���>+K�x6.{Q����f�����h~�m�3�����G�xBK/ �U-�ş�����f��Tq1�g�3QL�.�� g�d�t�fx����9T�E:O�sI����|5%�(���s ������w�_<.J�W�դ����ܽ}<Pٚ��@��7�jס�Թ U���~�Rq�A,�h8�1��H���#mD�h�w�|��,���Ğ`vQ�+qp�0�����9UlE��w�+Ay۔o��Y.GҐҮ�<��rd����!���rà�_��S(_��s/�EtO�t�6���;h�RΚl�s(��i�;�(������`�p�4s�̤fN��>{��^<H~%��Y�mP����I�	ww.|ɀ��7O�im����}.a��qցՋy��Zͦ���]��5����X��7��3U1r.��M0�>��6�?�l��;iY�I�sˇ�D&�-b�TQ�K�Z؇ِ�R�������*C@w>0k4 + ��=H�NE��u�D���n	�aC�5[c�B�o������ _5�h�����4�� �����ַ61&�}�ubZc�c���7�*Ϙt�y��](v��S���]��8`��Ɔ������);��{e�]�ۨ��o�ή���P��X���uLX���wX*2���%��R%ԷB&�^��g�.6��73R�d��Ϋ�崌�B>�������4?g�R|�:�I��d���#��jr�]�1�rw����������}5~�O����ǣ�?Q�}u�5[�����c%�F\��m~o�v��sa� ��;���4�xP��B��$��s���N�n��<ˡi�����?M�������B�����_��أ��. �(�%m�p�p+z(u�;�%�s��ޯ�j�`�h�!��FX��%��ү�L�A�^H���)�6G��K�/�]������k��3�QC�4���j�����Ɂ�k�>s�׊�ͨ����9J�M��J}T�~��+u�귱F��w\IY%N����
q7��3���ZY�R���.__���0.��S���c�6�9vQ����I�ͪ����9��O�Dz7+�ū�Cr�`p���^."��/��|ݫݿ����3�W2����1���VM~�"�F^�CD�_EH�)PZa�u��3g[i�:Iqb����G�V]l��^�S��M����fFo$�,Ы��Tkc��ERJ�xT%dw�f)+�X҉Ţ��
����c%�S@�MZ�o@�G�
��CA�w|d�"��9Y%��i�8��؅J�N9�)�U�s;K��O*´��@���Pq'C�Tf=i5O3�-���gOZ6���51$s�S��7�~L����.�Rl#˧�Ű)��%�n7Xc ��S�3�`�*�t���V}ݝmjfs��}�����������fw�Q�Io���Ԕ�@8�DxD~;��T����>���ԩ�R*�m.��ta����E��ӽI��1}�k%��a��U�5+������P�d\��1���:����ȹ�0�33Lg&6�gG�-kdV�H.W�dyN�Z:�=� {�o`���{�������SJ?A��=b����v��%�f���R]�6Gx��������!k�x:nۇ���m�G�5���S7�}j�[֝X%i����5VaZ�tq�ѡ�qVf.���k��D���X�u#���:!�;e��^u��e��aK�9�/���DP�=[���f�"<���Ain��|���
Q�C����Z�E�z�cT���	Q�e�� �ش��A�K�N�0FK�5����_7��l+:7��Cf���@3�)d΃}��;�}+jn5uPq���|�.Kb�PJ��Ѳ��{C�	���H�����#Cco��/�'(g�A�+�[�x� ����IvŢ��+ B]c�����SiR����v4`�o�4^|dG� J�sڇ�F3����{']�` �e=��6K����31����DD{�J.W��x�\��7M<��Pm�؇��.(n�g�{,��qc
�P,B�X7Ν�r9� kɯ>�A���Z�L�L�B	/��X�����/��s�� ��dZs=�xk���kp򆬴�]� }��+��.�4�U[�H���l�ɗ��w�o�F7n�7�S�#���&l���m��n-�A���GK0% *'�B��,V���kQ?h� �*y�xe�'�9dU@��`����іc�u��4֠\2�B�Yz�d��D5��&4qFN�?4���W�/ TDc�s~O%(]���/<s��g��s܍�ϯeY?��A�m5w��mjv/~����������۞��^��Të�4*�� \�!�-\+��
+�D��ӎ�\m!���;Z<C�7�XE��
��>2Րj�R,�k��{����4�����W(���yT�t��o�O�y�Pd'��jʙͯq�Bʟ3���$�N���Ln`�����z�\���:����!������
Ъ���t~Z�LC0��S�c�L��x�l�]��/��EY��j4�	 "�6�H
�.Q�v��+��i�����>��*#�N�o�,B^�c�����kJ����d5�+��ٲl`J�)�s�[�B6��� =��I�����0�%�(fD�78������[�|�D�n�I�n<Ӿ�J�Gr��9Fx�V.�֥��4�iV�3�m���;/F��l�T������ޯ<�<н����bΖ^��O\=� W��#¶�<�~h灶�д�	�%�Y�!J>�6o17�}�#\&Z��������L�m$�Y��ޠ���,�|��8���y�{���0u��H,=��C�Z��rd֪�P�0���q\e��4�V���L:���D���q����a�=�d�+�wPe%*��� ��	yd�SY{8�.4͚��e0�����1�h)�aR��T�A�~m� 3e��\�B#�k� ���,�6J�������Aw�t��ܽ�F��t��_��	����(���S�@�`���x�F��;'m���9��8� �������<\�+0��h/m���Y7kd!����q??<j��*�8ooG���iq��G�wq�6n��o����Ʈ�MM�(��c������:)���<�9/'�h�oTx�\��a�<������M�6s���^�jT�b�v�� ��Eƌ~�Jͷ����&��}Ѹ���$}�g]T2�$�\��X��X�^.;��"ۓoZ�k����~b��6u�h�(P��t�MjL�޲�Tr ��'E����'�o&�Λ��<���*V\����Z������%�sR���B�J!�Hs+����lQ��$LxCC����鱁<�*��%���%󚫨:������$α�T��v4�
�w����7M|���\v}X���f����Yk�[%�����̋K$�̮���,�7%��|�i�]0�ĔE�	�]"�O���� )H	[��"���1�����,��ڭ�{,=�/�V��@��j��qZ�ES� �h����P�o^��K��Ф�`���3L���$+!�`�zn���Xy8��3��/�.\|Q� .�`B���؂ǲ�h��vg^q�,�
��NB����`n��jB��KÙ9���w��&�o�����y鏣4���0�Ax ���J��UT
؍7tU�U{&�>����L^�gT�R(L��G�D5}�s 3���B��8L�)
	$VQ�僋�'k�Ǳ���qoƽ��]d؁�].����ۊ4W8t�h�����o�^m>�x�x�Q�� ���$��U��{R�?�_Ĺ}��v[��Ջi;�j �Nq9�,� ��|�Y~�t�o��H�:��'�wj�Ԅt�N�ЉS�hW��nwUݕڣ�2w�ˢ$n��y��7%�yb�B�#�/쩏-_���H6���)2��L���ӛ^J"E{����c��N����}Q�~W	b|,E�rʥ���yV.-GLg�:ߍ��� \��'�K��bN���:D�?�#����J�y+CP��}���0x��M��|����ZYf��Q�9�g]�K����5�%=0mT�J Зh�MX�'<�(OM���sEq܆�5��A�<���F�
�9���c��>gg�r|�Va���G�)T.���J�����q`"�^�3��1��B��+ԽI��z@g6	�(�$�_a���_��EұU�W}��n�����z]��~@e�T�)`�c���A�������2��V��&����3f��8r�X���D&nW0���{����7P��i S Ţ�A</�x�r�(lо.v��Q��1�X~)l�}�]t��0�9�������o1��z`�#�UJD∞�G�sܞF���}���6�$%�FM�{M`7���M<h91RQޡ��^�x�&�}v)�{a�����o�*�t�ڭ�f�eՈs�!}�b Cɷ�#����yq��{�����L�!Ȅ@�q) ���p����bL�;V�vj)�9��I����<
v���R���r�^�m;=3|�iG���
���z �	Y�n ZԈ�׌�p1|�*	�cf hH°���W���!y�]j6���H���t�1�ٖCѧ*R�Il�\������@�Jb�Sz�}Fvi��0h��%�{��g9��>�F!�@K���;��0�:4J3����g�n$	8�zNrgg"���p��kDL�1
�W/Z��r@����նy����1M���Dr��၊j˯a����g����Ή����y�X�������8���_�>̆�!����LA��8U�"��x�0�I#km�\ެ��bmq@��s'3T$��%�R-���\W�Ǖ�O�>+�y%��i�>.�רǊ��RN4��8���c����!�`~>�bL�VS�P)"�Rl�s%&�;O!@cN1��^����n�쥪���=ңL������6�@j��EV���iLζ�7���`�f���b��F%\�'K\ a7Ka�a�S�˪˴�%_�&i3^�CM��"�,.�eB�"�$��.$�KEQcYv!���l��	��+`M1H���\TK�T�X"�W"|�=v����硳��F�� �Pe�=��	0h����p�Nإ*�I�!q#�}r2:�*bD���l�$�M�gm���l�*?��|E46�-�FMz=8[L�8��Ǌ]���=�|���԰�W�Āb��aI����I�!�s�EI{��=vP���mZy�qϓ�?fBsRq�z�������l��ی�$�,)VҬ_� �%5���xv�,
���_c�w�ߙF0��#2.��=�B��P~r �]�C\�nc=����F�i���+�gt�j��I�BхH�Nm�ar��*�i,�]������l���m�q"���P��QTrl���u�}�W:Q��p�O��j�l�=2�~ⒹqN�OY;�Y��sBA� U�8���X�����{+9 �!U&0W�$���jº��>s"(r �*�Ϣ�}������z[�I�4����9V�`=�ʋ��� &_J��#�>A�s�g�_Η��|ZҞ8���?$��h���:G\~���劀&�ǬQ3qЍ��r�����Z�4葛��,wr����HR�H����/q�#%�fjpmR�/�qկ�w�Ը��B8�ܨw��V{Mi�s�����<�qVi-�'	8 z��WhRuM�<B6>��S�/�ޱ>��{��X"�4��\������m�X!�����W\�h���8>T�S�]��N��jU��A+��gI=9b���`���� s[��$V�22�q�b�j�!�K�4'vI�:��$g�f�-}������������rC�ZIy6CD�_��!�M��+o�h����pS������c�~���u!AI 7~��qgԌ��|�ZQ��{��h��`aQ��Vn �vtUM��%|*ṁ��xTa��yۇ��c{��n_��m���*��|�ˋ-���8�#aU"��8���[G���ʫ�H�Hb�@�0
h��V?xyt�����7'���yV����M6��'ٗb�"A8䱝k�Y��m����=��#�?�
���&�ib�7W���y^�x�oB}{�g	l? ��v�u��R�"������V��/�7�К��긶�i���7JYf@�_�h�jt��Y�!�N�3�yŊ����>L����p놞]�6���,�M�fLI8��<r��L������{�J@�z��	�ޟq��r£��0=',���Q���w��{��!{������Ҵ"��4�VȺ���6�� ������J�Q�"߼U7@�B�����TK�Q�<��r۰��Iě��m��]�|]#�������J��)U����!ocծ��?�f�p^A���$,�~���w$�$�d����?(#=D&r�(\P<��'0�6�n���H��+��>�T'jV�w�ʅG%���R�Y�:�T.���t�9Np+�W|T���ͯ! �������Ӥ��>����G�����D|�!&r�M��1�������h�ix��fI�m۔[��Ak�����=ێF>�d�\#-jn�#m�
��A�����x��f�G����L��Z�/�I�֟��m���V����zH_p�8��ŕ\��h��Bޒ��auj)K��2%X@^�y�1b���9:a��<2�9�ʹ�[eTI�C� ���ߗqHj鎚ǧ��Ԏ@픋ʝ�/$?�k�</jՄ�ў�=L	���-s�# 3t+S�Z`
���P�;�z��]{��`��>�]�C��o�SkM��ʪBc0����ޠ顃G$��o߳~�o����w>:��zՉZ�<��b������ �iu%5����#�7	%�L����v�YV
�L�Zφ����o�^�%"���vۯ���=�lQ�?e���~���EhQ���On���i:��c��7[�ֲ��}?W���so���M����N	Of(M��H�>��1{a�sRc�z'��ZY]8�����psέ�Ѷ@�6)���}��-j܏<�0�gF4���Aгϗ�giU1�ӕ��~팼Ⲯ�X�#�r1� - �(f���%�����+�AL�f���r?ᣊv�&=���.ZMe���踂(N�qG���[ۏU�i�Ko���04wǇ��l��	���'k�~�@-�N�䓬u� W3�-+�Ɇ����mV���a}���.+c'f=&�gZI�����������Sh��O�bv���q&��R���!�@A�.4LE�=@��'�ҥ<޳�! w��mr|�I�Cց�6��-F\�.5t�?��k���S)��v!\�0�_$�����D��CaM���&�P<������YmD�t��Xl��0��s������ڠ1r�
��	�|f0��,�JI11a1���|�6i��׌���-�?Y��@���w�?&�n���e��9�EOvr��K��x30��r��+�E�/\��ê�g͛���{�NcA66�,��2'����|pŉ��߿�\����q�h�sx�"�`|����PcC���	��0�* �(���_���pi��M�;fAө���n�(�M�rrm[5���d��
���e`�R����(Ů(�a������=��6\�mt\[K�W^�R��{�8b�B9}���5�/��Dm�^^˟�(����w����17ڎ��>���C	��b� _�<�o�Q�����?��f���x�Ƚ�f�?�b7d��`�� 7ê��hp/�/����OQ�e��9��ɂ�`]���ܙ�t�ǃ�Zzy�-��h�̕��&`��1�|�K7ש�Y$�	�#�����z�SHYg�d�Q���X��ط�r�7��E����x���9v�**G�?��v/�� F,���z�ӏ��Qa��NG��Rqi0��rw�T�Ȃu�o-
-x��%_��䒁�*��5�6N�vh�H �(�G!�nh�}@�D�2TQ�7���Z��̚)a@����qB��3�J���Y�v��Lfd���3)����x�Z��%=V���b��>���:�U����	��I�&c渙��#��mg񃆂:(P��*��`K Y�Pە�����/9�;Q�����哉�wQ���|�����$[p�ߗ��k�u� ���E샑l�gv>'�1|��u��F���l�-J��1��)��0�ra��c�6�nZ]���W��qw1�Zo�e�D㑯�����ݴ�P�������Ir7�V-�±ۭo��V�c��*����� �$,�j��D�����lC�
�1f��|l�%������E%���Xh^)�+�M��7�e�?\�hxpD��t�w	u���D��7�dwgַ�Þ#�w�'�'U`ۛ5S�\�<6��kn��Č��� �{�J��{��L���0Fp$^��K@�r�����6>���$&@r6լO�D�+\=x'Dd��h�y�}�X�v��a&@y��3�k����fe���X�|0�$�H�ĆhN��d�����٤'
��s�GvZq�N��E�K���1�9	^�g��f�ͦ�� �7,(@4�'�ڬ(Rrx"��A�S&0wM���+i�۰���*�1n��9��x^���@�$i�"��Lf#�T}��}����`	��EvN=�A���d;������a��%߉��w~w9�b�#/2 ����L�e�1��� )ɐȠ�KSb<��
# ���t�;
�\$�,8����X����?B��]뷦5u,>7�r��h� |�:2�������,בf{'((LY�Sh�VJj&�:�zxY/�&>���PE�����Q=LyC��Dփ̈}��G2e)Ћ�ǧ�����҅aإ�
PKZ߹����:wv�����hg>�F��B��|;���?���G��JIh��9nNzE.H�:��x��Wg��Ȉ�D�j��o�+�|*1�ejaLKb���z��d�=�u�[�
k x�d"�	�Ҧ*벍-�,yv�h���<� D��m�'�AT,�-�;�
�2��YK��ݐ���c" ��w,�RN��?o��}K��Jz��o3�}�~��A:NN��.[�8ι��k0*x��!c�̭�(���t>@�nDCͅT�A����^�*s�H[i���(�stʸ�|x��c�S�(p}��#��r�0��D�O�}+{a�������78��ι�6��FV������ᓞB}����-xI밽������Y�#��H����g�KT�>����{�3�_]G�R�)E}z��T��P���~�@E��-Bc��"U���80R���ێ ����Q��(B�l�r��Ys�rj}��l�@3�M����ڲ?��dߠFZ'�bo�zW# [�P�r���"uڤ�$�w3�Rm�zBU�|
(�G��|�`Ke�Jj�q*1~�`3�O ��͇�}�1e�ƻ����;����2�	��<lsSy�t���gD�!p�{Q�:K�0w��}�b��%p���S vt.ǧpZ�x�*05s��Q�����ky��P��e��b�o۴*�^@�b�o�D�͚vi�g�æS���Hל�c�D�Ŝz<"���)';��[=�h�&�##z6)��B�'G���M;���-1���?�p��,)�IO�-�R`$7N����vA@�'2V�J�����wm��c,zW�>�5!�tN^�e	���)>�Z�.�,d�����%O�zB�Ӣ~~Bv��2��� ���<���6����A�E�B8\��ۘ�{=g`�?�NeР��Ctڥz� �k���� ��#G���(�N��
�������	�R�,Ԗ��FN�yx8a�(��M��G�{-qIͰ:�9�k���-��7;׿���Lr�r�U�o�V�u�u2F���˱�̒Q�g�:Z����J����HًC���M��ܻ��J�Þ�2A ��K�e�Vι�ۃ�G�iq{#,7��'��Tm=ҩA�vT��[�+���r��z��6�X3�A��+@+�b/M6L\�rb��)r���1������n I������8t%������|��b�!�S�.��8����O�֔���ۋ��g�G!Ԣ��|���K���Y�;���V� ]ɧ�gsqڱ����w�&��f�;���v�
�i�@����;�nZV�$�|e�%*=�Yp��}΄�5�VU���A�̄M�1g�4�����&���ػ��[�|����L7��Q6�qJ��V����V�B�H��/s� �����k�+�̛�J���j��e���V!���{�3�j�?:��Fz-����`Կ�{�Lk'7nR���"?�2�jr�BD�Q�=x�Rq�-��&ނ�)����a;�5���5rsH:l����6r��sG����N��c���Q�CH�m���ҍ����UGR�B�"9ڡ�TbJ�F4t�&�I��_�!��w�Dνh�e܈F>d�t�X�����:�C�?:6����H�ѱ_�ќ�?���	�[lmW�\qU�������y��Q�(vS��������kAu�ZD���P�+�U���%�
�����u3�"����3����VOi������z;��w;8�n��PD�|м��Xe�Z��*�L��nH�c��G2�'U�k}]Ss�l�?D�WA�1���vtg?F!����������&d�z		��-���N�u1:��W|��R�Pf@U�r����7��|��:LКz����ĭ�G�>4
Gk��24w��㻏Њ�r˙�OWWV�g)dQ���5��fI�U0��eъq&A�M�,������
m�}Aߢ�O�1�bplMǷݐ��(J�K�g]�nh����oJQKQW�4�_-����m_f̷�U��\�?�a�(խ��?	#AX���ƊP��<ܾk!�3˽��.�������^T���Yb��^O|�l�H�(�P�z� q�Bヵ��>{��b�וu�
!�bp*�}�{��}��͘x��u��Z�8h�)5Ƀ��mǌ��wq[$�YLٶك����b!o{�L�V4 Z�����!^�� ���ο���t
�G�B0�k_H4ǩ�B'Xo�D�.����B��>�Ѷ��]�����^��bM�i���P�~�>��Tx�!\Ġ�3ϣ�#��~�N�Z�!�����vG���|�
@k}��9sQpf�6I��~���p6|_��xr�Z^�-��&ow� ���XO�J�0��>l����!�%����X���W�H�8���M#�L��0�>5~�QJ���X�?�&(I�Ĥ�&�E�hn\$����m�� =��#�w��2������]��?M�k+�Tc��r׏z�n�.�.j�_I�ګ,H*@O�$u{׮��P�2&�tv�mM��1oyZ������S~w�_���)�Knh`����Ե�E�'���vs4�Ы�
e���2;�=�	�*Y��K��@;�%��(����'�s�A��G(��ҙ��<��������cpvt�����D�`�r�y"Rp������n��w�q����5Ff'�{e�D�K��kσ�b���s�:	>��)ͣ�|h��`9��M�dD`���1���>�z�~�G��c*sAh�3�ڳ%�W���zZ.�p�$��,�>"�S#|������	��ʹ�~']�
��*q�:Ps�����nb��q���l����1[娲����,_��i����*�.�*D�������.�~6H��4Ԟ$���m�bv�	�1�:�D)@������o��#�Me���̜'���]�u�B�#�:3L�oY���y?]�eܤ~����|<��Ě*��.O�)*�`|�L]�ilߤ��G��w��
f�m6�.���Ϡ�i�L�B[�ą}x�����=T��q�Pڅ_758��ѵ���\TG]�P��OvG��G�}B�����m�敜A�^�Y�D��f��H��ŷzĻU2ZZ�opr�
W>�f"��_fJ9�yA,�22)U��d~��P@T�Ѭ<75�944�zk.m��*�{�_��#B@�!�������2n!pܟ�1P!�r?"��}��A�G�
��P�������WN���K���`���Ʉ�,����d��]0�l� e��Sp{�U�l�t�����֗Т���#-!)4B2X@D���;���QM@���	U
'�P�����A����{�X`��첸:��',�4/�*E�W��nAy������(���x�W�wy"�x�T4]�q���3����Ϳj����oF�w�:� ��_� �N��V��5��Q��@f��w�if2��JpgG�s|�V3J�e����Q�� ��Dۃt� �Zm���%	���<�y�����+n���Ǎ��ݸ�M���CHĞO2,�CT�}nzD�'9��?��өr��%����x��b֘���-u�rMm�??�ޑu����T,f�\�G�7�9��u�G�J?s4���шw�?�0�\S2Mh��ɽ��+U��y �hP=�da����/fp@Z��[����m�z�Z��}�"�}�vn�e�����K�A�&U�*Z��B!��������������U�Q����.���0�N,�H7��Δ�nb�����g�{��N����t"���9�٘��4nJs���P�Ca:Vʵ(�3�����I9M�R �]F{vO"�^�35�6��'Ŀ�_�ĔH"����'���*�=hS3}�R<E��M��`�,�U/y����Aq�k��=�iJ�D�����N$�#s����Bn��3��"3���D�*:}�>��~��5\���m6��DS�r<(��̤a{���vN�����m��"\O� j��t����`�I������!u��P����ч9ZT����֥gI2���d�����J|w��B���~O{ {e>���D�J��~J�,�t�%9��%��{1��)Ur�i���������SE쟖}I��@�/G��f��|��ꤨby�28�
3%�<F��5vW_����#׍�믇�Yh7*�Ґ�6i�vk3�TS�+ZH:���]ա�u�}�g&�����v��£g��!]�T��?�	�d@0��,σ���sP1~��S}(��v�>|E�3��e�Z%_��
ML�>���#�� h�7����;��V���$�`^jj
�S^�� Buc���4�h��L�����d�p��yW�I���C��,&�u�|�s��XP|���N�v�
y���x)4��8�HV�?=�8�r�I�	]�3�=Fe���
��X��ty�K;������g7�Ŀ�	�,����b}����Zճ�`�s�����B�+��8CV�yc{�B�`2�y�]!N��m���(���(>�!�mw�mg���m0{/�F�0�^>���RZ`T�0�g�a�ȗ�1|�eG���7��~���&!���!xM�T�oU�L�K��(c��!N���I��!xᐾN��'!���~T���Z�S�����9��"���$��@�{/�M�2U_o���(��0�����oP]��#�h��Ѱ���|�>��(�Ԁ�^e����Ty�F�6���a�뜰 Q_�Mi�՝��G�Ξ���Q:�,+cs��0q�AZ�WJ����1+@�L�!.�a/���/�,���	](�%��;ں��]���[f,7�{9�K0�'�a��{l���eA��WD!?7h�W��A e�d8v?m̔`��ū�>�*�H�[O?e����5�b��Yc��9���6b��VGi�c�5�3:���Бx--5��T	��P�%��Q��D�'����ǋo�R����&�y�������M�K7��T�\n����$�"f�`��z����
!rG�&{�������yNx�^�	EV���%�#օ��+69�V�?_��"lD�܆�>.�TUq��!M��ֿ3SE7����6)�W�Q_�J��I�Z�a���m3�yA�jm4���-or�j��5��a�!W��S2��!{k��/�+��&C����_ �[[� r��H�q�Y^��⇚\-��]z�GPG��gj+�Fs�:=��?b�x�e������.�4pb��ؽ�+m�g8�&U���Lp&�K.h_9B6��4r�F���!1v�(��ָ܀��f��#�8rc��b����Pb�L�r+��,����:���g|�"����Bk�^$G���f�+��TͿ�8"�����l�<F9g��gb��blm��
W'����"��3��D��R��M{)�I��4��~��}��j�|*뻋��&}-p�hW�/�|�󃦪2�5&f���ѾRx��N��L�X���Bl�Aݣ�<�����b���Z��C�o!�s���K�'�v���'5(�O#�q[`>�֛�p�}�E:�ǟ�����}ٜq��p�{J7����*��+�&���=��� �l�w�~�zK��+1wg�RM�k$y���-�[t�D
���n���b�Ĵ©��Ke���������N׻J���!C�[��ל�$��$GfB~��dҠCj�
»9ae�eᘜf�����`�����{�;̯й��K�dHf,��6�:8�Mc��'�.��}@�p�Q((�>o!3ɇbC�uIǚ�,1��P�!�W\q�� �rD�h�F�#;�z��%-�pM3T�B�u����*ᦃƿ�񫅢"C�F�=���#���oȸä�.n��34'�~�Į�ʕ�M��c��D�}�Y�TP���MCj�?�P޼�W�pOm�[��nYp��(�xj����ү�m�`�%V��k.�a���WgF��tI�{c��>4��!�[��Z��b��Cٸ���,�ͦ���[�q{��	!�YLGXQM�E���;Zk�������i�P�ag �m���w�������O��a�Q��׸�խ4�ұ��$k�_a�7�!����Qp�f� �L��/�:��@���m�����-��s�'q3�B��4vx�Ъ�ۂ؏EEDtH��&\��I[�&`��!��w�����B��F�0*4Ab�&���
o����5=ś�.������!(��d��k�mpH�,��AD�d4��(ϟ�AD*�A̟a�4`�<��
tA`��	��
�����i��"�}>���Vȱ��St�'���1Õx�����
n1�`S�\�zDă�Lv����'X�/::��bq�4l�C@|� �Y�}>� �aݮg�K�bZDK��Ӥ�G6҉��D�t~yU[���`��<�r��i"<��<%�U�[LU��(���U��M)�:ǎ{�q��dgYb�;T����Ё��L�^�p8ˆ.���C��m`go-}jڶq�Y=�P��WL�����u!���q.Hlީ|�߾l`�}G�$^2�<������Q\ T"�O�l6c��d�g�n�/S� o|��w:/��R[�w�x,�n���2'��~�gwu]�׈u�s��!��0r���x�y~/��ma�~�zgp�_�/�G��Vc�Lv_DH
ޔ�ܠ*�o���{9K�:` 0~��Ι�:���C�b�
��NC.����ͭ��] a2��@՜�_�����E���VNɩ�9�9Ɛ:�hv0wɜ�`C	��٥O����߆����
4�8���zi��s�[�ZUM�/�w�ZSk��g ��:�aU>��7�BA�R�V��I*��D��4�P��'�^s�+���9/i��22���P���@�{j�ѝr������쩮$�aE
BSe���p��H�	�ݢA�h����&��P�a�7&�v�N�u^��ڶ�h׶�8��]���t>�����`n]�����(��-xǧ��)����X^P.�;�x}��98�6��(��P~(]�O)��>��\C�	�Ή��$�$M@pf�Q0�Tby��� �>��O�J�}���_��N��ݥk�#�o���L��@�x����]@�I
+uA0p�?�BGh^Z�����`�%%N�q�s��b��Hl�ߍ��㱑��"EX�cۍ���;����h�}"��Uq�j m>�D&�:��C�U�JOI��DZ��3P9<����]���$��z��VB�%D#_�e�}�	����-�1U/V��K[s���]�D$��������~�Ք�tݑX�׹CyTU+z���#�OI YY�S���*��/S)�~�Ō]��Yx�uݥ/IR0~�p���=T-:Sǫ����|u=Z}�H	q8������\x��mk'�"�/u��d���N�*� �/ ��f�
�!i{G��?��,W�Y@(o)�����{O��NX[�U��q�F�9��;�P+;0CN����ܔ�l�4]��c��l~�T-/���%Ga>И��R@�ϓ��G�ڲ�7}H����G�S��������Ը{	*�a��c����6:�ˤ�2Y��X~�Fi�����p�%PF_V�p/�:dv����3�X�0,tS�-Z�'�� ���z������ުl ��o��G\efr;4 s)uN�7�V�^&���)�f�(�E���w����$l���@���\�9ag�'�`��6}^�ktm�b:�2"b@z�v%���^m���n�b1�χ_g|rd��@;�ږ�O+��BY��A�~�|���ps h��'T&����in�s�%���5����5��b{�o�BET�M�!9��p��JH�'�e�P�~ca>�8%��+2T�*��> �xkh6���A%ʘ�j�LhX��RQ �� �N"E��+pLpg�W�̅B0��33�EϹ�s(�����8�k�N���Ջ� ���b����Ц!��F�>?-�˻�D~q3|�'7����^8��&�O��q+��
/IߎětjS�§���G��G� �y�{ZV8W�zA�=}�̋��8�pI��UC�dߘS�	�?a�w��.���}_��1��������YD0��jԆ���/��5k�t�^;5�;�<�)���4(���!�'hZ �=����c�b��c�����3Q�_��\�V����y-=l���;�#D��0BJ�tRfq��A@G����U��O�E�{b\VO��:��?:-�<�S�ԹƲo�f>)-ɊJ��Z-��j*vL7 C#��mF~G�E�6Q/�8��(�WsP���\�* ��+f��������#�����.�����OK����(���͹�9���:;vj�c�T5���]BD�w%�`�u�3��.d��k\h�_Zg����n��QSo.�X #n��X����0Ѭ����%��J����Pox2�j��(��:���B���[�rB�2�O�/uQ�ø-��5�gV���݃
�S ��x�p��K�Vw�d{���x�C�@��J(Q\�PwuR�xAp��O�P֥��k����/e�����&l��睆�V�������v{������	���'?�w}9��4Q��N|�%[��+.Y��������^)P�x����@�Syd_�p�P	&R��sa��}{i�+K�0a�I�5m�V-{Y�s�`�/ݠ����h�R��;&�TɢPW)���,�[�Ւ�<P�6b�\��: k�ؓ�"�ϖ X��t��GG>�X�xy�(a>��`}��f���e\��r)�+>�}_mi`4+>����0ck����m��u-�H�`Ӫ��ַ;
�~#؂�WG0����U��ń0ɇ�'٨3W7۵l������,Vc�yb��"f�Zf!C�X�</r�A×�))wA�f����PDk�#zXN� �p����!��g��S�84�S�p	y]5���ф�XlBn����>���3[��
e���K����λ�:� �rд+E�D��B>("DUH��u3������F�����5��������J��߲v�k�m,ְt�*k��Ѩ�5#�<��?:g�x���%�7�*!����b�H��u5чK#�����et����"�J4�FTZ��%Y����*ĖB�^$�E��)D����<�(�h ��7�pMK�OC`-Xf��O��BLG�ɸc��Fz����t,�5��4ԕ��x8%��;�ʀ)�%�7l���+���7΋Bԥ1n�Q݌e&R:�e8��$SUδ�J�����^ؚ�,$jV�p6���3�� ]Aޚ���>�kG����1ݠ7�uֆ����w����[��?��	9X�i4ʳU�<	)馺��뙹��&�?�z�!8\�~-K���mZ���:�@,M��kg�Kd�	�՝`��].W% )gX\��-��{�(v��5�a�}���}�S�Mbcdh�����K^��/d�jY�Z��(�`rb����ǃD��C���fV�H?��n�h.j����t��>Д��#\�fj��l��HPWUO��yH���,y�L9u�R��* �� W;r�yW�@��/��O�'���=��vӀ��p�E��5�pz��p�"��Q(3�xA�V�M;+�.?Q	�l���+;0Ea`-����p����w�tYP���9�G��i����MIǥ7���=A`�9�죉��O��J�T��ύr��C�
�Ա!J��S�%Q�,XR�5> @�~�w���T��p���+ooCjr���[������{f�0���q�l�r��L
��Ip����A�@�s �A�� �e�����.�.��b��&�̷?�_�+)7T���R>�o�S�:K�:����Tά�t-Y*lt���kDܺ�8��[	=���� ��~�Ր�j��mr6��<�>��qb�ď��|a�O��-o^�өNmVӬR�j�U#PğP:��f�0;����z��񇅟44�I�.�]9�E�]3o�Q}�p�	&6�K��y�Lȶx�Ĩ�d���~�(a�#>�ɉR��p!���,�O-ò�*P���-�KX����(��~+�fH���Bg�(?Rr�+yv�_�%�fF:	-.��y'��Y���dj쉳҈:㞀pfzZ9�>�ɝ�|�#�&ܺB�v�1�YU���r��1��H��ډ��3�;�2�Y�S�Z&��d��K;��I�$��yR���k㠊X��+�d�,�5������`pB��&��G�lㆻ��������2� �U�YƉ@�^YO�J�������tY�RCfbt��S
�E6��9 x�v���T:���Uݷ���H�!�"����7��օ�4=sPS���ZK�����1*JW�!@(�>�͹�9��O��>�Xq�]���!��V�����-枀��!�+�͜�rJ@��ID���P�
 _b1���3AqQA�Ք8��6#���2A%�t�/��s�x.2%�wJ���GH.d$а������-���W�!��G`�.?j�Λ%?*I9Fū�	����)�m�$x5=I�o.l����j���3�RO�_GR����ϼ?m6��[Ǜ������J9x��$�T��s2�0"��m�0��O�;$_�@�`a��o�S�����{,�J�m����ɉAЬ�����]>�+v�!Z �����н�w=��(P�C�Æ����~���4��A�/p��I��`�s�`�lF�V��(�,���ᑋ4uA�Vf���5�t��`ʵ�N5{���)�Иb=!8;�/��q��d)������jޜ0����+�����B��(D��b0~�X�U��Z�y#N�Z�=�~1��G=WP��gu��_P|����I[?t���[Iz�������aX�J��t�'���s���:L�9w̤��
�Y��u�~W1w�#�P�{i'a�Pu��ؿ?�+����y�q��~N8�_����X�����BL��Ͻw�Yۙ/(�A�t���1ýK���i
�B�lM�+J<~��3)I��b\� *3,o�t�y��(��U⭵@��:wX3}7�ю'���2�OS1=��%��@�%XN���,L���r<����h��LdƯ���U�<WCg��x6��� B��3��4a�xk�9dN�W�?�"q��-i/�A*�rT#��(�r�����%/���6k������Is0)�`�B�+w�f�������G.��#.T=������ ���ǉ�^v6�x��O�=�.�ޏ��]~��o�����}d
\5��$�#-�=Q_x�(t�]�1�;�'7�K�� ݊���7���y��mL
�F���H��5 ��}G�^��_9�V5کgf|+;�8��
�xY���L*��V���*I��#q�/�`m��q�DV7Ә0k�]T�0�[,��`��#��G�� ��:�æ�qN���q��p���IK�.g�2����v�-��K������6��	ߦ�@�!r(0�$nljǚ7	��*9�H�읅�t(xf���x[���c��=)�V&���T�~&j[{�/̏nA�ĭ��M��	{���א�ɧ��q.[��J���@���I��ƀ;��Z�4][���0������F�7��4���j�Du��8�#�~hM�iR�/�$h�'�e^0\����,�>�h���a7jc�N�a��G\}4k����F_�;��K����3͹MG��	�MS���hN��0E�vԾj=o,jLr�L��;�zXD`g)����TcA~�ƛ�[�V�����gʥ%%�z�(��R�R��ձ�^�:>�i��\1Z�u�e��FĴ*�lh�Gq��|��i�h�MJ^�iszl���i=ly�L�+�x9F,���J�g'%��g']��>w�Ey7��y=.J�(��y�ҥճn5�o7��D�U�`�|!���CR�K�vPD��\l��S�2b$�-{>�	7`�t��*C�nT���n�=���7F�����̬��8�%;|�P`6?X��IF���d���l��l�?G�ޠ]�'(���΀�@ 3�o���lOJ;F���{� �A���H"h	<~J�Bn����������{�?R0�{29NЍ��Y$��j���:���T�����%X�C�5O� ���9��:���n�ny�K�8%I%}�lQe3JTh21��۞��$
5�`������:��嗃4z^��S��ġ�n�:K�/���[w�u�sܝG}��?��-�c�ξ�"������N:SzքB���rC[ k쉊�'���ٚ�ѵ3g�]�/�8�I�>�M�Π�g�X�;O��)���G��0u��K{�֯���~ؗ�F������q��9�dk�Ԟ�΁2u�2��1���Q]�i�F��(n�;nv����������T��6j�Q"�V��%x�Γ�+�@�U�TZn���Z{����{�����
y�8��$�=��+7?T��H<��cv������d��c%p���E�9�ʨ��t�Z��Q:���G�fHZ���]����� �u<��{Z�̯���V�l��9�L����ޕj�'���������Q���^$פ�̠G_
;d`F�Ӧ��0�����F��'�e�lD/oR2��*�
`�q@3BD�h���5Ջ��M<<�O��#/��'�������[�߮�YZ$_�h�4��.?���k�Q��$�	�CQ�/ C>�ăo��s���=��[Z��Q�׬+(_��� )�
oa�4"�q�%�蕽B�+l�h��y�����E���7��w��s�w���a5*��T=#J��V�9�5���.T�1���F
�=�XH!_�?��%�O@�E�O-�P�'��6�|f�Ys�FQH�7��#6��a3g�Z,��8�� �o�X�������`�G4��2��8�z��Y��̜�:�2d#�	����F����C�(���}MU��	�H�^;�?�`���D�X���Z8��$,��dyX2��NPЁT�������)_'�d��?Ӑ.��]�jqc\.% K+�W]�^��	3`)=y����'aPt'�4A�A�۞���-WF�V;�#�W�1�H=R�k�'ʁe�G��;���\��.�΁p����Q�Hf#ޠ{v�G�:qՕ�	0��L.9F:����-|�����v�ׯAI׸�Y�%�a�H��9FD��M����=!��d�2����� �7�d/��7۠���W��Bp}HI�*!��@��}��"��A8�%i L�J�G/�A�)�}��ϲ�]�$���N��[�����]�-bZ� �k1��Q������=W���Ro8u&��O;
�x(�7�i��U�
�a=��z|�լ�3�D�1����.��5�i�~��p���s6>¨��IH}����1��u�(vJK��P�b�"�gҐ����F�=�8#���7���Zh�uN����NE�����Ȝ�p�[��3yܼ�ԬJyeT��{	h�
.7�3�1'�{q~�4���V�O1}9�SJLsG3;��4���� M=��(���_�"�G,��-�[��n�n
kbHw�7<3��c�������㜾�D�'/
�ʵe�qn$ ���n=1��㗮�8���U�d%�X�R2��FL��ȓ�"ٗ��|�����O���q�z��Vˬ��%�=����pד��=�qf��8M�Mb��#J�x�Z@�7-�jkQ����{����������a����`��������J���_Z�U,PQ �D��*�`�*�Ƣ��6{���[�m��i���G.Tx�2��C�SҀ\<%f�^/\y�7��i�,VL���yK�%��Z]��	/��ͦ�3�&"��]��Q.��|y��
���{��;d�����H�|��O���2s9}LFQ0�V�	�	�=9��(���������Z�}؛�K}?��@�����0XH�Ď�d/��c#�KVs~N���2�ɚ��l,b���.�R���<�GS�F�^�,@����&��ؚ�x����6����M�b{7�l�l��8�rB�C1�ф���.`�@�oEw�V~f�bg~U�>�"7�kI��AC>iE�1�2c(���>N�5�wƤ��E�8]��j�d_�Hb�&�����Yx��WVٻ��YE��#����B([�"�$���U�̮���4�]~b@���D&[ࡺ�V��3-4H�j|)��e,􎺞��ht��UEY�.�y��s���˴������I�*7�8�☆A���f9��z����-M��R_�au5�K(�O`�#֝��T�]�A��w�#�<3=&Τ�Q%�(�����~&r����;���Z�A8�:4]���i��xh��˒�Δ�W�h��aƺ�ͻz����Z�#:e����2�f�vJyƍ�G{1ӑy�i��A��WD�X�h5�5�aTs�o�)����*�@��O9����c]���.�	���K��S�z�b$Sy��-쎕W�pk6c���*�I���|޼�%c����;.���a3
�t(�OF�]���0��Es���4X��Hy�jo�G������kΑe*08h���S�&C�-�ݩH5~�NA��A�@g������S[���W�EӈT�:�M�Ci�)?�~����6[B螈��z��F�w�����=��O�z7>NCK.V�l��9�6a�횪���b�;<�p�C�?����#.a�2/`8�t)af�m��9��gc����-�_�*Dzv��y8G�����%r�>T �z	BI�;Ȟ�1�����w�D���%����=�;F��n��H�����">pY���j�A:C�D��syNY�ٛ�?m�"S�ۑ���h�e�@I����*YS"�2]C��xʛhRȭ0W���Ut�)"��|1=A!�i� ���ԕ�¼8w� )ϺZ��qZ���s� _�1%��<�&h�S�sC��it��qa�L�W�Z��E$؎��L�D�A����m���c�,����4�?5"5>�� 0�ƬC���bVgQ�#H(��z|V��ES���i2�E�j��?H�N�!���t9��;z�S��� ��n��K�����p۾?��
�fB�R��ؕ!�&���Ap�T}�}`������+��6�Q\�$�v���:&t�/��P�Fh�mGh�:|�����I$��.�Ka�
=�j.�IƮw"��WE�)|�����9�}G���"hｃ5�?���j�@wI�DIS���
9�2��*��6'��]�x���r e�E�?��1"E�P��(��	@Ķ�ط�Aq�;�O<��C"���ar��j�I��I>I$�(oQ�h��������`���� ..���Q�����1D&#'.E������¬�	����G�+G������w	/?�x9��ّ�6����I#>y	C�JSFO���{bڀ��yM��tJ��3?�]�/9�u���+���Á�;�u|��&�U��W�5�>1�T@b�U���ɫv"�� ����n��g���L�O_�Tb=���"��(�d�´듒�<=��J,|/����j&{�b�m�,0�ɍ�0{  Xmq�mh0YX��������"0dV�k�}ҍ��Y����mWh]bD
�cN�an��+�V'���l�:�(���nj=8�����h��j2x�.BϦlo�#� %�i�Z�'�W��
�V��=� �U�eKZ@�ndT�3r�I������:g8��a�.�8܃��'&ޚr����x��w�Z�L"�hN"�6w��N폅��'�{R�ѱ����a��\[�����9�D噷Q���#h:�)zC�9Q�qz0g^! ���\mC�¥B��镎����_~�X//V6B1�4��_���#�z?םT�5V������J~�h!�+��;���	ȋ��>ڿJQ+���J�a��3)�-���)�:�9�w'�Y�&�_���<�-)���e�ҹ�_��dEvB�+N�ׁ���l��X x��q�6��nt;�%���<7Z��">�}����X4/���r� ��k=�~i!�ذ�c>{6��Ү��� A�@�4Æ�b�-��s��R�н�Z_��(�����id��zt0MCjyNjW��"�N�� ����H��ȜC���]��<�����
�5O6��R|���w�V��ಀ�ɓj;����|D� l��t{�$���;�ޚ~NSv#�ީ֞5q<@��צ�Z�I
�<�;����Q0���j�f����C���S��\��O ���L�R�7�<�ʫ*�!�*hށ���
�6Z[=;�:~��<�3�(y��`9�{_=$�:�����o����v���I�3��.�%A8��lLs�d�V<�0��� 4:t�c�B�Z&_ՠa�'$q���U��-��a\Dp�V`�ڍu�bÓ�Tg�T�����:U´^&��Q^�2��Ryu��$D饉y���D��Dŏ4�uj`����~�[��50idjn�YM'�8�gR�j_.��t I�r���+���#U����I���/��Kڿ'ߨ]���$���q�x�A��N�D1 �Qw�tW�By"�����~���V���ѫ�j_d�����K������"�%l#YCld(33x��cV�����N5�p���ۺ���|P�7�B5`���'�jW( #{��C9>��A��Zm#��ҽ)p�M�s�����@��t�?��d<	bFX��a���˃6�R�ԡ���Y)f�?�H�҈�hl�|�a�����ʱ�% u2v��^��T��*�_s>�t�c0�@�|9oJ�*�4E8�a������+�M��zyJ [�jA�u[��0"�QxA�G�%2���x
\䨻9�ؽNʥ�k�qxY	�z��3��i'2��O�{���~1�ug>��Q����'R�`S ��Ѝw�&���x�k�P/�O���yt��f^t��$�j7�먷s�3�/G8.i`��tT���^�$~,7=.ӆNֈ�0�	ڿ���d'J/�ގ�<:AW>@�����kN24�V9>I����U�Gf���%=�h��dY�	��cq����Vn3ڑx�\ޯ́2N�_�殺zg����|�����k�H" ��X��3pW�Ε��4u�w��$&̚�����4�u�S���ؽM�ܯ��11�ǃ��$ ��M����R�(X�ڨ8�g�τT�VC� ��|�+X�ObB��! `E,�f�ZϽ�,s����7&v-������qAR��s#�L�ٌ��b� _���f��Y�Qs�Q���ZP�P���}f�N5~(c򑦋C14��D#q
o8�hc��I��Q�Y4�!�p�l����׹�|�&5ro�$+@�bDIn��[�f�hd_=$2��ֶ5��XB�A�ނ-=�Yx�'/B��P�=9x��bRa�]ԡ1KC��#�Z��$�f��j����s�+4��|��o��[�y������><����&�Y��I�i���o��5
ȷc�9�Nn �Z��aY�m�i�čC!��<%��C�D,.����fN�hF��d��Jr��9䭧[�G����Z��G>Đ4	���N1���0`[ x�S��e��X�e`��0`L;�o�b���oa�-���̦U��`jD�g��ى����)A�%:��������p����E�@9r�;��GO�g���(���?ZD�l�#��Ӣ��i-��E�y�TX�J.�t���i�D�5
ʣ� �M���0�%����U31�eܝb^�����s� �l?{7�*-������w{g;,������)]�/g��ؒ�����Ō��ފ�F'��] �q�A���n��.�_m{��uI���tR���a���;~����Ogk�7R��Z��x,�	�M�~�{C!����=���N����4Fy1�|u����/�b꽋B5�G���n^C� �gVc�<wHnk)rP2h6҄�=��b1{��p��;}�^yd���)�_�sNA{gRU�_U��~����=�J�d��/�)��2n�Ge�E�F�(��Y��աnA�XS�i����x#ތ;#��I��P�;H���N�	D	5�ۍ�,�J��tz櫪����W�N����
��Kc���u����9��Ql�^x���P����$������$��B�X��~=�mw7{���L9j��z��{
sdJ�ٯ�������K�Z*_A-����D�T3���ZX������h`���6�R�������	-��y<��z���0�V�±*c4Z+g&�����T5,��MTXp���3���O�� ��;��c5.�g;�,����C�� �bY_��E�v��l���+B�#뷆ӆxA�y���u���lM(��I��0�T�/�̟�#�0*���K�*�����`"1鏍.j��:K���A�utܐ,����'��^���o�R\I&�$6S� 5��������ElZ�$�I��{���A���9^�}���qe˯<�}<��IX�.��K�kN�Sr�
�uF�֎~�W��$Q�Fش�Vx�4�H�}�D���L�(���N�I2흓�Z5P�~7^�B\o1�\��o��YU@�Cn�k3bk�;h��2�m�tx���~KT�ޘ�0���N|���L�Y����ڿ�y�'�$j?��������y���c�����9�i�x�u%�-�ڠ]Ǭwe�T��Z�Ј3�6��q3173s�8�T6΁Z��2O7�X��x��ܗ��鉚J�ub�2_v����k�[�����ڸ<��{K.'ss��z�f�����0��W-����n]�
2<��w�,q5��2�U��(l��Dv)��Lu���"fd@��`Q$��i��ֵNj�L�%�r�
����T� �=L���`�pB�XQ��5���91������-�?��ɽ��)U��ك���,��'�4ʞ���ه�]]�d�O9�囦���1��u���� B�N\1�x�N�&b`���,tDJ��#�o��\
:�Y��W�K�����s��Fl�\�.�m��vG[Z�k?��o�bC���v��͐ƫh�x������Dp��^�q�DMS=&j�J(!	�WC��f�]%�f_
k���%xu��~� ��O#/>wB�˛��WhZ�xt�����@WE��~�*pBZ�+*�.aQ�k��ǖ"���0N
N}�c����?9���v!��>:0j hOb�M�E�c�9������;8X�K��_\�J�S%0mѵS�do&��4�s�Ng#[�R�qO������a�%��6SՆ�E�[��,�l����#�F�N�b�ܮ�hW�AEu���%-����K �����i��ǩJB��`�P�� ܀�$AF�����<� ��fhg�Y�b��]��������'�ͦڍ4�5�~�Ta�I�<"�ߴ,�6����3�����pm�"�6�m���+8>����B��<A:�6�9~:�G|���)sd���8��ga-�c
�yח��g��8x��qɕ2M�r���s/�:�w�~h�@e���T��=OϒD1a�^)��#p_����s�!m��D��Z�Ϩ�2"�Я^��%0���2�����7? h%)���u���l��F���_C9� S������Rd�9I}f��ntսM��.������_�t��m ��$	�%8c�i��7_0'�x蹈{_�PK�7ȣܞ�~�ib��%�(D��3����F�g7ėP)���1A�0���X�g���jOZ�����kT�t�ܭ^�J��FI;N�]�U��.e�B���3n��?�����C�=����=̯p�����6�u�Q՗��+0������9J�s&�U|Ij�Ru��-�8�E��~C�Q�0� �U�T&�;��W�a
w#�[FOT�*|�m\��̝E�����g�'�En?ܴ?>�++թ)i5���3��q�Z�ʯ<�UQ6g��Z��EM�&��@?�M�b�o��&8��g3�F=�e��y4���;���|R���ڮ6V7��Q�U�^Z?> ����r��-�V���F���,s2��@ �1_y�k'b����%� ��y�%�!��Ѳ������Y�O��S~�7���w��P�εZ]��7U��'Z�q��g��3�Pm�����ه�MXIR�g�s�	�\��J�h��v�VT_2�#�xWM`Ngp��?�d��_�q�^C�&3�:��jX�#uIĚ윇AGvX:��5>�s�:]$��ƥ���'���(���)�"`Ue7em���$_��Q����O��&���g-ᓊ6(@a�e��ߑ�t��K2�)��&Բ��y�ۛ����-N�	��N��wW&;�W��q��Һ4�ѯs���H�-��A��=��@`�a���Z�o�E�baĔ��b�Gl�8�ڣ�&��W��jT�(��P�dg/��ef����0�2�~�Rۥҡ���$f��+�T+�"C�ˤ���p�$��CO�R��!�����|�<�C+�H4�PZ��W��=�S$͋@�~�"C�R���Vb.��>�P����p+Z�!Q̽��긒���&�t� �-�9��>�P8dzI��&��iԡ%(�&�g�(.3���EO�M��EKDBW=u�%_��`_z8u.��ۺSx��L�����w ��.�<u�S7�Kx��	�o^�1k!������2��|ס\��@D��qkhBHd�i�iG3��e�1lw�=p�prd����Kȿ�9R��B�!��|��ip>1�L�&���XV��&_V]I��y3q/0�����1��&���tG���2�')�\��]�l�O'�O����oي0�Wjm�{ʱ@�e0|b6�t�=^;;\���}^�F���x�f���j0���gw'�_'��j�lMB�:�kϘ�j���V�҆��{��R;I�����%��y
X­}n�|��b�ŗ���p�?�QMu;*n¥FW�Y�������F�ɷ5�N�΂N�0��L��0��˿ 8��-}�-���ԍ<;>0)�H�E�Af�if�;�����- 5�a�V���n���Ix�*l����M���p��٢�s)�-eږ���\8�&��$���,�k��'�ù]I�-����k�fG����`�\rI��$�^�\h��[�>��"���H�1:l���~j��"�pSF;��ϊ��=l6녅k����[�晬 v�5�W(	���5�#c���6tiX+���;h���m��λ��5	7A1e�v?�@]0�l�8ԛ�vV꧗�\mp�����h?�+W��0��W�d�=��ON��&I�|��j�"ʑCy��I)*H?��DG��,^��uNv��.*Tpg�ހ�2{�)h,S�n�@�q��R�b9ٮ���s��IiG�X{�{��D{-�)u�
l���k���b"O�`X�:֩YY�e6A(ơqV�
��ge6tf�6<>L�(�s��_3���z��[���=k>70� �)��SX9��g@��)L|3Q�(n)��3ӧ*�]�N��(U��jLiY%�w�έp���������ˎ8K�7�~ųBup�L'��jJ��H�at�d9H۞�0���� !@��;�"�� �K�n�����E!o�<�K&���A����~���Nh�yl=�[�u64У������[���Q�h�(���N�J����(�����H�����>�+��������#��(��]f���W���%*{�T>�"�!s�Q�k�F5`�"������ge2d���"���7���ɢr�M��+=����$u�b8�ɻ~*������������ `'��m���� ifH�揎��ǧ+�'f��/�9��nS�xȬ����u˵�e�}��H
�,�R�X6)����4Ṩ0":�Zl6~e�LM��4Gq�(�Rp�^����=@�����Ho��@�7���Q��%��7yl(�*mQ<Z�κs������|��p�'�K��!���&N����yѼ�Y�%�����u��[؛^��)��~�_V��lb;I��FN+��;�zKV	�E�<V�[�Qt�v��|�<�}R�����k��E;I��ׅ���X��#�$\0U9�[�6����q!��!����ԍ.�Rfp�X��eC�ݷNimo��,�Mi��_��N7pĝ���È�O����	ķsܴ�nuߣt����#�' E�G�bar{ҵ\���^5�|^��Z��:M���;w��Xd��Ga��P_����*���+5����ٽ�Fe��<4u��o>�%���.pw6l<G�51anxZiI�q���l{�zGe7�^F(��sUV��9a �`j��jx�	^:�s�+8����
NiG��I�t:����{a�ԫ��e�X\h��������ճ`ɉm�dm1�d�J"�1�:^����C���� ;�Q�"9B��H;�dgڨ�41L�7��E��ºs�^�cp_n�W��3î:&`};��)�Љ����1���!)�9�ɝ�.�q�M5��#2%�2�iH���E7%Uu��
��WKn#]�y^�,e�<2!I�8G��yN⊣"�0��l�x@��&��g��BM�z���3h���ϻ$��y���Ք|!�R�c�Ӕ��4�e��fDr�����b�Y���|���L �{~P��������2TƐ�3�ȴ�i�[��6�� 򶂝�:�b�c�NFu�i��д�kz�!d5�)q+�-�,��	�k��T��18���f�eq�}�I��k��U1�NM8�20�#}^�	⹬d��*��ʴE~)�{��s6\`��7�GC�	�����'�6H4eF�(���k�j�k��9%Q�o��X��f�f���AN��0ޢ���c��a�؏��kr�(�����&r�"�i�r�VENYcl�{���.�ce+���FGƥ�������(��m�X�����ix�dw������^�U�-��`��`ŝ|��X���6��~[�g�v!:D�I_��l��G�S�#�/��8CK�'7�#����Z8|���"ufΛ������y��ڀ��
���+��{Mo�,�� ��L_یO?=2�Q���mr{?�\���*#�hV��?��t�H��whh+
�P�"c�m�L�3?�S�-���W��ݏ����K1���bGĦ��� �/@��q����ch��r���^&�ۜ�!���a��Z/%�:0�@Gl�p,+�h�_�������.��a��f_�z���ƨl�L�r��HQ�E ��<j��kM�l�P��e���$p�g��Wu�Y��F���X������TC?j���M&������#p�@�2��h�0֒���B#���J�3�/)�o��y�fS%>��iė����Q�|_P���D^��3~ �|aٶz�d���}�%ۑ�v�T5�c��*��Ô0�i2���cN`W+�����3�d����<�R���2Q1>�����Ώ��hJfD����L�XZ�z�
.:!|�}�/J%/-k����*��WEs����YLQ���):I�|fO!�|�����/��q7�m�C��fĒ&k��VH0�9����E5�OL�r�f�V��Ӓ�!̫���4�h�شTX��'��U^ ��ЛK����:S���͝��a���LJk�����	��T)���Ъ�>�q�X�-3>��R�y9����|�j���ܧ$q�?ҹG�d��������Sa��{���|�=o%����d��t���f��EkL�3E�s�*��5�A��������� hg���Fi�=<P�]�TU�p��@�{�)4N�Na=%a8��ʈB��e���\�O�B���&�E$Ϭ~
����Wp����T'����J�P�b��C_����kK�����;��	m�� lt���=ǂ�)b�=6��H�X���i�@آc�&�ꗂ��?g'�Z����N#.rp!6�\���;�бi�hé:J��b���>��&�Okw(��9���]an!�:��������&!��e�ff�FA� =UZ1�
��g��l�/��ߣ��ۚA�A����	������_���Ԫ�n��գ�HDC��w|3p�Oe��7V�e/���Αֶ����j�)ԋ�#�tm`��L����f �B��'�*��e�[R�V�[ت�k�ό|/�]J�i��?/��vt����e�+��:u ���L�A�}�r����M�t�Dy�#XO�� 
=����iiGA(aA�/6b�0�v���-�4;������c��ē��a%#|Y7���0rv��(sB	U��L@�P��c��t�S�8����	O`�7��$5���k�OtLWk��|]���(�]����⨌����B��&!��h:)����d�c���fj�pfI�]�߬�5s4��w��b#��-����p�t��M'ir�)KA @�,��3#M�!Ǹ[�_��Ip��#!��*J�@tM���!�x�@�0z���x!5��S.����^,�6�NQ�'6#		�q24[yS$M���2�s/M�չx��h	����������%J��x`�b�'�[�����K@���0@F���l�B�����z�v%W)&��Ɍ#5���=�����}Z�s���:'a3�U*sۡ�@�u�?)}��6m�]E�wRjk4���h���0��kE���}G����҆�*	�HCR�X���Ɯ��2Wpj�$i�zſ�Zx��th�[���BI��uЁS�h�˹����S��� �+��ܖ4�N��L��+�t�I^M/j�jE����m�z��F�y��1��j� p�*#��Ѩ4��u���w��pHW�_掟#��J�iz���F�լ�ڀف�G���oRd���#s�����n#�O��d(��ȫ�Ob�ǩ�;S*$8�����ғ1x���t�Iy?�䕸+fv'�Q��z<�����8��!;��L�F���O8v�wxwE:�V���
�q����C	�����2JI�B<��9OM�WC���C"�"����Tv3(|b�7�A	iL[Q�K�|�3G���l��������JI��,-Q�����i]��lc�=����d�6w��P�󲛘���)κ��V��q!�wМԽ�p.�u�%�w����p	�',o,�$�p_G�w7��h�6S�isi���m�u\�Qg�+��Q�b����	o<S6z��F[��I�6��8D9����֣����:�w,7�B�P�D�����v~��1���yq�gM۠:�_y�������T2~%��.��a.k����`�ę���+��T���#����r�\�
,j�H;�~Ts���}Bw� 6�q_:�z!	�O���qn�M�H��r����6���bԝ٬6C�S�=,�$t��!��c�jF|�:�`�(&�{:U�^�����F�z,'�Xz$�n*�(yK{��b�l.S8���J~��?��/�����hd4"Wg~uŖ�p�>���\b�2�.��մ�n�'es���	�<����$�'��l�(�L�9N�I�|A������Q�P��|k,J4��p1U}�͐��a�"����0���_�ff�����h�Vɶ=��7'p��ʍ�0L���'B��>-4�պ#P�]��jr9u����v�S�4�,������+�,�[ċ5#T�Ḍ����i;�
r���u����qGW�B��'8I-X���6��������7S�ʉ�'����y�G*W���>������3I����l{ ��u\3�I��r�%l:��ۂ����MN�64�� �.�9-�C)�Lo���ul�08�7�u�q��e�ɂt�'lL>`$���5�_�R�!�]̬��\��H����F�p�uB6,A4O�	��*Y��U�3|J,�z�Q�6<?ro�}�L��_!����/�M�n�ܪ�b��m�>=T�z�\������s��둎C��`��0Q+�zz�h'	4��,�x=��}���@�m�r����8�x��n-v��:7
�Y��*���?׮��%	7�m�:��}��o=0#�@s�9,�x=噗V���4��.!�Ӄ��ر��g{��U-E�4�S���Ti���9k�e�|W�a� V��{�B2�,�r��,�{�O�������e�f,-�qn���"u���M)�z%�������T0��Z��l'2��]�@b��|to��R�}�:�c�#^�8�vb���]OSٺ6z���
���V�ҿ���<�V�P����}�VCY,J -P�T5~K��s�8r��¼V��s8�{� ��۷S!�r�M�-���bv�!H�c�Z�A�t�N?��a�C�$C7�q_4���7!��xE�$�a6���'L���G���:��mV@��-J��2w.�:uNG��x��v�m6:���T�$��(ly�j��bTND��mL:6_,Xj�ϖ�p��]�0����Ȝ��m���<A@�,��+NIşq��	E3��	0���']�A�T�Mh�K��sJ��PM��k82�=��y�O���5p�X��kV-��i�_ִ�G&O�]�w����\6b����ZO}�}_��~��h��.���#�٩&��]��w�t�M	����E͊�'�����2|^���G���<�q;R��A����#�ܤ�o�.�)�1hQ��]� ���l���D�/<Җ���~��'�逓���j��	́��n�f{[R/������=	��� �7���$�9�w��TJ����c?�@�G�eR��sn*'�{�A�����Q�b�O�9����9L�w���B*�}���w�skn�8������+<�3�1f�-OAL��,vo��5���y��O����z�px�fp���Bצ�2��m�T�56Y5��H�3�ЊM��-H�hy������ɬ�Yͥ��/"rY�nZ��E"���Ӎ�P`�(?")��\x�d��`.���Àa��>�&�s�N�E�l$i�Ͳ�}8Y�9,�ij������ɟ��qa0��]����(ST�OV�����y�.m1ϼEE���Gq��>�%��hn^_�ն�ԝ}y����)o����<�br,k+�ӧ�Vc g9,{��"����~}���w��5:�����_��Y��/�?T"9����|�C����V]?��7�Qs��ȶ]�A�� C�������J�h��rc!��V���*�9��������0���}�T���I���W�D1 "���t2�L�5�(��f��w��Yy��Y�/I��w:o���D	��W'�+�_v↲7u���d/�j�$�U�:|t��^��k��9ڄ��S��������Y-�U���+A?�}����WɡĮ�3e��'�iys��v������B��]"
��*���uZy��H;d�/����	���Oa��ۀ2PJ�~C��?�����x�
	�����$@-�����V�]�g�h���+�����}��1qWޔ��z�]�V��[�5�y_�^���4�^'�5}��cہ��xI"yXӆ�����ͤ:��N�5�����b��V���x��2��'W=kSM��1ӧ����fvtd��� ���Ѷb���D&t��Z���b�J�)%=���(f&?�	v� �z�L���@3l9���7=)x�V�Ϳ�AUlP����h����(uj�$הݥ��G����JX�Ĳ� /[oxt��W3�D棻H�t����_�,���a˲E�ykU8o���H5�i�ه<�s�����׻e�Ǖ%]U�����;�7��p���W$YZ��݋_�9�ڻ?��$���β}�P�Ha~R���9��P�7��/�e�S!�߬5#�O�vu�6����)��v����Yj"ڸ����V�ZawJg�o�4+�}�#6�׈e c��"d�-�w�����[� @]cѻ���,�@�w�ޮ��S��b4k����}Y���}=9�����	�,�ژa�o�:6��ՓU9��o���e��}���ҭ��F����tY�����V?����Z �/2�X\
^Q����l����[�k�_0����L��u5��$�-A�A�VJ�PƊ������avstc��g?{K�Y����) �N�[JZ�U�=��%t|ʈpLc@yf��G6���f����\��|%���ץ]o�c������D�?ꓸ�N���$^.��:�Mw���A$T׵��8�؀uá�g/�ϊ@N%Vc"��=�!�
�RV�f�a��6k`i^��'�T�5��s��ٴf���n��L�cn�[���D~5J(���Τ`��I�r�lj����U�l<&w�l�T�V����HY�ba���B�G�4�n �s�2��턎�:�E�a'Gx���3��\b�!DL�m3����M��t9bGXZ��<9yN�dU��l�~zی�"��b*_@x'�z�η2�]��l�=Z��6�7��U�Fo�b��]/��Kq�� �jj�4�hGӑ�z�[�H[^�b����k��זА��=�UL���2�]V�ύk�2�Bs���W�����5L��`�7�%�ܟi$�i11�1�aks�g_pg� ��<��D�I�
"�6#�+.Ыu�$�!�ꊋ� ��4qAo.z<&�� "��V��Ӈs�#�yn�Ҳ���2�nr�S�>?˙�n�N/\@�P^V|p�O���<)�ߜ�}M{ӫ���R��-����j��g�*΋Ĕ�\r�\�j('c!J�z
�v��:9r`_����lR?�-��<
1�$#h�p��?�XQ��D�c��U��b��߻aC��Cע*/��$�S�4���,a�oɻ/�|�^���u=ЌM���;�o�8���1c�'�s���ALʾf��l#N"����MY{Y��LF^\'v���}���loy�/8�e�"�D�1(m˻�
 �"ZЂZ&~,�����������	aF���e��i-�j�&�П��-�(��up�J]���v&����|��Z������4\D7�`q,1���̀�0�^���g��*e��2�ĸS����jt���4E�����JqV�k�:�����){�):HC}�J�d�,"7!�M��{�P���P����h���Z-�(�	�`Gd��p�8->��)�9�aE�8iU�L��g��{G��z}ـ�� ���"�A��hU�U@|�ӂ~,��
Y�� �沀&y��7|����X\ĕ�Af"����+N��a}���V��`����x`��o�꠱֣0�VB�y��1�:M��P(�\[�tM'�'��A�:�_6��ؽ��G��ջ?O�+�ڻ'���T�O��۷Ytơ������V�GBצ#q�ƘB
���?��җ�}���覑ԫ̰�)�F" �#K.���uZ