��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cТ�L �~!�w}�O�ﵔ'��E�L�i��=/�/lq!�.B)�Z��Y��sP��CYvS����+a_o�&��6�K�b�
�d^ɮ��$z�U�*a��4hb �'X,+_(��
ԛJ�	&z,��������uzH���!��Y�<��+��w^J�4P�5�'Xa��h���m�������^oi��G�-7�/G���~Z��~E>;�wX�d�*\�n}�;�iph@[0s��!c#�6���a��sҴ��PW�w�Y8�jS6�O$�u��>�¼䟂&4=�^?3��1�Bx}�d��{��Ai��b$b�F����������I��Y��*BĢ��:T�|}��uT�V���U����2q��L/��2�B�Y�hq���9�z���	�Q��A:3r��I�F���[���#i�vE� �ZC���ES)Z!�q}���o���%�Fp�Ȓ<X�Ad=�T�y>�7�q��,�Z$�����z��^t����_�0����Q'5�w�s+���j��[ҭm]m�d������
�0��bڷO�)�Ŋ;���?#����dㅿ-�<�ﾏ�䯊�L����X���d#�N:+�n`�������kzg>!�v�0�۳޹��%�I�y�&H4�)pqIp2����9�5�L	�TB���U_X�$"��MU�u,���R	g��r���Xw�F���yy���JA�if�@��·!��z��__(T�n`u�D/|���E&�xZl�J�(\<���P�s�!�Χ֥��ۯ(����٢,���D(4sdm�x6�/��k���BJ��R3���P3?[eG��7������s"���y#ֈ9�BE�V�!N�9���ؼw�����SV�Ta�Y��>���f.�v�Q�\���6w��P@Ok�&��mY�b�X����4�͛Y��d���2�$�S-�KhG-矗�U���5D��7�Ŀ�Z9��g��Q�[�-�P�s��Xc����/*r�*�7�F����h
�D��uF�+��g	�k��h<� ozp� �7�LvW{�Oe���E1�������_OWɬs������^� CF�w�z��f�o�AYl^J���=�W
�R1_��4��x�$�\I�ty{E �h�V4.���p	Du���K�*�Qź��mzF���,�W#G�o.�.��*�,�ּ�YаZ(�]��Gr�Eo3�jz. ��#D]�u���[�D��	��2ei�;� �J�nX�{hr*�� ym�b��zS����N�b�m�?� ���l�@?n�K*�,ֿ+��kSzN�{�N�֮o��H��YF>�)��l(-�6\v��%�6 �1w�D�.E.��W�M�lo˩\�u��NB��m��H�i0S	�����h0�W`{���쭠'��V�Iy����t;�T�[�|d.(~�cGd�����69$/=d�n2����)������֨,q�e�󝈊���}��F|�2�[�'��ş.fy~�&\����~W� 6�ԙ{���֏���=9�,�'y���:�?=me�$0�,w����U�5=�Ǳ6ϑ\�'�J��!��|�}އ�Ib��t���i#�ơ�.h(��?�����������!=m~��5!0]Ah��=/��{h��ʛ��s�BCm�.p+K��(;
j�Y+�m���{t��1?\Y���D�5(�P�]�x;������R)/���g,��i�ع��F
���-atAZ�$i���Zٚ	����۲�9��T�����ڔ�c�"���ˌ�D�`-�gjpN	^�*�*27�U��Ț�2��{�/k��@ŻE����*t���Ə>GHӏT�U6��;� �R�7�Z���a��Lό:'x����8ẄmqJr�r"Ԕg_���ZƸ��ǀ�I���)���}��[�0{��N傰�>�w����GFn�	6�5���z֞��J
�e\ ���#���`~��*u�
dٺ�|�{T��7�F[]���&�X\���S�:�J^�[���`��l���(��T�uET�Xg����������y�l���9��R �����-�h6L@W��O�Չ�E9����-"-4���� J�rCx�r�����)m�p���!2�ӳ\���i��U�Fp]�,�%�)�O��Cߕ���������8�B�6m���<�I���'�����y�DHLȕ��@�Ԟ�@K�H�$6�z���Y���j�r��ƚǢ�b�]��oå�v�ds��=@�����O�'%疑���|<*�w�k͋#��B�`���	��~곔cY��3s����^D�����Nbde�R�Q~Vq:�F��h����6G|t���^b�p�'���]�.��@�D����T����D��* d�췷7L��"0Q-��ĺ1�U��j�NaU>r��x����)���ҕ�����B��ϒ.%�m9V��?Wt�����|C�N�e��D��������p���+��&V��(N����%�ް�K��*JL4pFlr����x��%�r�"Il�JP&C�)�Ŀ�ַ��I�m?3릕��Kk�3H1e���PP�4���jAJ�'љ�!�u�a:�8����f��������{ƛ���mq_V�+�ڣ������9�Qd �K���PT4��sv�Xg����ߡ��H��<��3��\`�+Ɲ���BmkY���u"� �4�A0c�",�A���q�%'Z�155dc+���'��T����|<����- ��7��۵_����r'�g�����w�p����q��>;6#�����P��	,v�Z�;�k7W�g��P*H����a��ӌp��6�$����em<��Iוּ(}N�?:�=���%x�M��QP ����PAm�[�y(�>b�u���x��3�[�R|�I���/����z�]χ��8��eȂ6,ƃV��1�S�rɬH �d~,� �̜h#B^R/�
��+��撠AI?�%/�����wk!v$C�)�8Zװ��S�bxb�.C;# r��%�(g'K��!��Y��JF2�����z���E����޾�Z�k�<�F�+��ZdK\f��|�x�<���i��?���1K��,��� ��?&5 �?�K�oWe���pBJ
b��lы�.��;�֨/�Ӟ�Qz
j�|�ָ!e��?�=�L�D��~M��|P���zi) ��T�+mi����YN��W'��q��_٢	^��׌G��_'�?u����^�r��|��!#8��y��;�����)! ���M�Kw�&��i~����%D�9�PS��p��)N�X1�;uAS���~q��P��>\�;��~�"�>�]L�%��L��i��3q�z�?^�곡Y �DU�1_��h/wj���i�b���S43�Db�t�aY^VlO���$Y��Z�S���&�x�X�6�bK��>����0��`w�lj�>��_�'A�h2_Y��!���fĄ�� RCoX�tKW�H���b#��ck����JP�o�Ȕ�qx�x��f*/�Q d�:_I�',�p�7���+�[`��nށ燆�綈w�:>�2�@as�{��_��5�ݪ^1�/)sg�i��"���a���ev�ۂ�t�,%���R^��Ĕ>��B��kh�EG[!_�-���g�����M�m���݊�4-׃�sz�Ǌ���\��q��׊�����k��]-�s�5��rw�ĥV(�~��&�!m,+i�,Pa�.$��)t >J��pP���C��� �M�YFA��0��Y?�#����hPT�O$\�kpR�u��5��-]��$N��s��Q���R��O��S9o��М���s�:��t����P�9�j���c4~�CjK�,���pb��a����e�<	3���f�㒨�Kc��N8bB"t�ۓ�����'������Nw�G�	�8(X�g3��3#��p��^v��!n�ۦ��A.ni�a�y�黆���z8���r�M�D�,����A�h�;6��fJ��9n�"�'�q�&�@\�LpK�S����(�0�����3;N�_�pg�^�|��D�]�.��q*��ۍ���qd g�)�+��s��-�F<�,��^�W�b��X�Ʃ.��=:q�i,���##w���I(�X�t�����.����������H����d6�����s�
߉�����<?��ޗ�j�sԡ�Z�����,�	�$e/?�o�k�`�6$c���6�罫�TX��5��Y��f#���E��NRe�%�xu����|D	���Zy�]>>+}�ǂ�D	Zl6W�eXT��U�a�3Όu�	Q��0�\9QOf��e��?|�`邏ŵ�1q����;��-���䄈��DK�`�G�6 ��CWuU�buF?��wX'���6D$c��55o~N��r/�g��~v��y�9)6�Z^
+3���J��Xm�vr�Ew�Tl����]�'��<�-C����a~�-j�����3��e��,*a�c��L�mg�h3[���8��Hp��r�{���Tf��T�$�V\�%o����G�D�5)D�.$���ʚx�OΝ/�q&�-�����;��ez��o�#�B�p�H��םŲ�����w������:��ق6d�hG3V�`p�S) ���Y^��|ϑl�%ƳGƕ	ZZK�j�j�Ԧ�����N@���C�.�����yWi|w�/��_�A�Ww�浄�:�o���F��3�b�T�j3˜��8��X��tO�j�=`D^�*<l@Br�$w3��k��|d�S:��@���=oRE�O	f�
wy�cgg������e�D�e�����k7�@7��K���m��ٞ<"�JL��h_E�e�� ^r��V8ݝ�љ��n�(�h�������4� S�f�߹�~lj2-��s��Bc7��KS}�%I�N�\��_�63�R~�"=)��`��.�x^�{�6_�.C�k]��M~w��K�{�n ��.zȇ�gt�:6$��}l�P��D�Pt�y�S�;��i*��+agx�2�� /���\��y�� D�龊��%j"Vj�\�&f=<�:V�u������tI��'u��qYU�˕���/�1z�Z �1`�lW�ۯ@VA�{��R;����@{Σb;J�ŗ��
rk�
��A^�I{�`!g�x�φSZ��6Q(��~F^�؃vL��<C"%b����i��e�+A�� pg�NVP�n����������}�|�l,'����\�H�Kg�m���.��H���|+3:�2T�U��XdL+�t����u�T��y���X��Z����!�
qP�'�Q��w�&=�:�Hۑc�l���ഷH�åA�\M8hi᪚O�Ar����H߭�S@p3�����7�'��f �C�����[�uO�8w�V���q���
���
ܖL2��:��g�	ꞙ��X
��H�o�+L����­���6(e@w���3�r$�o� �u ��z;����f�Ghr��Rk�W����n���^i�ܚ�cL�?�Hű����\����Մ�������R*Ͽ�:k���l+u�+�%]�1�ي�'���t�`��
�*�w����2?�ӧ!q�;i�ʊ��O�g3���&�9v"|�
�	�� �e���8����8�s�ie��*�w�G�.W���v-I�Y����N����%s1z��CU��A��7u��<���7�P+�fss���JǷ��͎���f��ksjo����2T]�x�������8���d�֝� �קR�c6�!��hZ[��઄�/�!7�,بp1i���n�J�l(����h��9��䅸*ŉas�ҕ٪<�k�CO�f	d'u��jP?��n؂x��s`r����*����bln�I�¼��_�P����|1��bL�E���ذ���x����Զݫ�!����h�-�<�[+�h�L�^�і�@��O���͒]8����	QB�.��(�~�(c�+��$R�L: �g��ˤH���vwk*�9��+N��O�m��8~�<�qU��L^��J���)&i/9�������e��h�����#��ı���Pz˚�]���b����p%uY��eP�9Ed�UL�BQD)���*8Am���q���Re:׿��GJn	�}7Y;ŭ������i�ٸ�)Q��f�~7�}�h�V-���o��0чl%��8�4�g��&�V.�OP�C����jP<ȴ���_x�!/���dn�7;~�n��*|VhFeX1I!2�¢�`7� _�q�^j�ϣj�[|o�M.CtX.5n�"=��� �0�lmk�54�eKg�+�R=����t$Q�'`�R���]�?=�]�����q�e*�-�k���ς��I��ktL�z�{��寏����ռ����R)�~�f�jK�bq�G��s*����v2��I����.K�+�L�ޢ�������Df`�'J�2�lF��G�����>g��e��cB���[{�`����
��s�
@$<��R}&��~��>a��Es�Z	�i[�=�U/���#;��9J�RЁ��&ԓ����snA�R7m^1-��\kn����-O�ɂ��p�������_��-�j0Rƫ�[��K�w��K����� s	~�u��Gbѷw��6l�>�]Zb^�h��-_�=̔aK�|��W�X`f���eL4VBk���T竜l	7��3�����kd����ާع7�Ebd�m�X͒�'bw���U?u����}�%�,\ʺ��J�ڌ�\b\��!����yU�g*!��o�2���9�Dv牏al9�rR���p�H��F���kr�".n�ќ�'�u^�N���~�~��!-�z����~>�I*��c�xg%vM�B��,�ROĳ�\:���+�Q�)�w����k�����k���ڪPi�n*)+���gb�)���d�yf��rx;"�N��vf<f}��� }
��d K�ð����0#���͍:^Joj�*"�Sc�1�@7��5�l?�vgi^(j�Q{���^uǬ8[�����eଃ�8O��'7���yȏ��XBk3~l���������^�Ց*T]E'	����uY���$9����cps�ُ�(��ێaf,LZ��8q��K�L��;��=�8����x��rRt���1>m�@��xQc��"�n���с׫�����������:n ���]�D���sq�焮��j���n+�9q���M��&�f�@)�h�ר:�<+D�gȳ6��3is�
��kit�qǚ�ئKCBˬL>�t�A�1��(I�a�����ܺ�䨵��&��=RB�\�b\%$k�=|c&\�5Uv��+-O���&�=�����l�XI�������ت+R7����>*�������A(O�(���ja�e𻵢��E���1��ʬ�:���ii6�����3�V!�ז�8�qǲ`���=�]t:�5]�b<�L��Q_11 s�d��ӳ^[N�z/l�_�/���jK�es��0��,ķ��������F0h=�5�Rs�fj'���5�&б��օ�������1[kX3�}ă�OִE�fY@��@	�=���eE�t����CO�*:.� �6�F���S�		��7Äu�|ɴ(`����mE��	q�t�I�����\l�;���V��d�=��WN�(̴z���}�1�K������OE[���jˌ�?���t�Eŗ�1{[��@Ml�Z(?\�2$��u��gqβ>���K��#N�t�f-�/Wa�D=Ȣ-!��z�M����:F�;�xV�"�g���>�V���D�3��1By����G݀E���H�O�P�+���i/H�^�J^�8a@8st���6�>��"���h8����1_$D�|}Mo����K���Y�cג�F���{�$6�+��Y`��L�EFS�S��r��|���yL��r�J�Kl�]�4��Q���Yت��I��07����ɂz�l�'& �s�8'��p� U��	[Bi�<�+r>���?�i<(��ix"�҄,��w��߬�\�)+3/H��ma�P��*�P�	.����1u�B�Kɂ�.e�[��'e�������1�t9ac.�t��r#j�Y��E�.��L��˝��-^�?:GN�gi��X1Z��h����	Ə����6��x�����a�K�mfV�I<$��3J)�5e�419�rE�Զ�,���ɫl��LV��v�7A��f�Ż`.�-���̏A?g��D�K�oM�!��6���P��{�V-��}��P��'�VH�a�_�Jp��N�,��GQ~].2T�:�uPhE�������G���ؾx͜��`
�������1%/���bL�=������U����g���y/d	�J���-g�����vЊ��X�|yRG4�^G�;�ߨٵڸ��8�~j�ڇM	M��Z����{�GK�|$+��4p��h��ߥ̈~���mH��&�ʁ��x��%	��T����f�łϳ�o��	��B\���/Y��*���n����vC���Q��f:�z��#�޺C��~i��g�Ǜ1��%��](g�?Ү�����^��h�QF'k��.�͐wD���a�,�׭1�5ʣ�+��,����A4[�[b�H�ڰ���:��-�k<t?��7&�I@�_�ϭmO�6��X�f�j���u`T�{fF�+k+��#?�w�������i)El#�ʵ������9d�2A�(� ud
����Q�:����+L��>���B�*��ܡmZ�,��9��a��B1
e����9���rs�#j��,�1��kNSh1��� �Tj�8���G:�#�ɳ6��I(p݋!�����L��v<t�P���4�Vz�"�[���R�j]Brf�AT�!��T���פ�|�*���=9�;K��!��c��=����Fr����OV7�y�;�Q y���, C}���X]?��OƧ��^�p�R�c�FS`	�dU��Ѫ�{n�_m�Gڃ����0��JQV�����e�M�p���N0x-�e:r�h�&$<oy\z��ׯ��+ţ�Uj�4I#j�BZ�J��\�C��3g~~�z�����եƇwy�(�>2�7�?J�n�Ī?�(9um���6���&pu��fE����p�����p�2��'�;����vdXx����著P�v��X|�fP�����>����H;���ep
R6�W��JU�2b�����}�I,L)����LKK?18J?�s͖�m��˴.5e��7Q��R�)_�t��� A�Z��j��;��rf����i����7��t�Jk�
�f�ׂG�d�+a��>|L���.�X�0i(��-�vB_k��
�W��$y����Y�*��p�y������a���Ǡ#EW������0�����r*S�P��?G��e��bT�U!j	�����?r8��t�������k0<,\pn���u��\Q��Z��Z����QĒ�Jʉr��#�U�9hg�w>��"cX~n��H�*�.����\�������b� sA�E� ���?C!?�-��9��KG�7􇦃)�P����`��Ґ���)�=\FH�����#����=�7x;!�X�Fq#��ŇG$%�ɼ���Y%f�R[6�H�qmV�2uWz�9����n����!D����A�D���b�\-1��Vl#�[�=�����g������a_<.����ޕ����3Ns@t�픊��R�C5��|�j�}cw�M��r<v��va�b� m�.]�TV��D��=f[���%���Q��7�0Z��a'�y�zxd�0*G<N�ደ����nNm���Rt,�K5���R�;�Ǜ�Y��+s����i�eo�����3]�,�G�I�7�
1+��1b)�T-Fv]�	��MB_�x���k��L��R��\� 4�sw�����^Җ�r'}Г�grsb P{K)I�J��q~n�F��/���ٌ��	v)�}}��3���{�ֵJO�P��t�{��m �� ���#5�{��bv�M���ks�;�8�����$�흩s?�T�	�P-k���k�ā����u�e�؅�����*x�<F�%�p�QDp6�CӰ�s��W(�L�9O�-���~C�G�@f�wHd
���>����� ؼK*��7��G��;$�W�b�~�!n�YH0"�H�(�����Y#� ��y��( KK])rUh�2����W�-��v7U��iJӺ�cE�������x�U]S��<��Ul �G����%X8PIV�}���x�4/�N���C.��1�7lS0&~��GG�qiq@Z��ᓿ�<H�H���\� �0{30��n���AHu̗#�*mpl�D���_�O���=�~u�"��G_����1{�#��AN�s˦�Z��	�b�w;ɫ�������]�9�V��iX0}�*%�����/�1\[�����?�;��2V���ٝ��"2����!E��r���r�XX'�n�-�ϩ����E!�|b�w�XO�.+����@��s%|B�f1��^�r����I'i���J}Ęk�2�:�hi(F+�bH8b9��#��|���kD&�a��|{u\'{h���Ǧ�6}�3��ٝVۜ�T�!�."�A�м����ڂ��;��=ƣ����8x*�M_�܉v9���'�i��@X�ЇZ��>��λo�r�%��u�r�m��㬀)�@x���8Q5R����)�讒��D����Rm��kWޞ�pfu��t��cJe!�}m� �?b�R{�����ڍ�9bj��,�`�!����́�8��p�}�.�4�+s�e��c�I�D�SY,9�����.by"�Rk�w(���|�`�?6ʽgK�]*�Z��ss��u�˭���z�G�F<%ˤ��jفǻ=���{="<�ej닖��bئd��{o!g�&������ڤP���8�� �h������M훞�L���/S"���-uM�!
�LQ�eOlP�/�ScQ�ȡ6}m��Z�ܼ9��H؉������:���,�[��H���W�2(ci8���j���SR ���Ρ3�Y!��n��P��K�����b�54��\�?�n1����9tZc�\m��Ɏ3���Y^7W�{B̫b�@HcU��]���|�U���p����E���d�vE[F�!��A��F��-��<��|�*xa����o���ee���a�j��F�(w0�.J9LS>!��-|X+�d��{�eY������$t�D(O�1��Ł��O¡�u�$�K���9c�4�?I��%���ew���>	`Y��3�=�b�?܌�ƭe�ZZ�	F��F4���0�p1p5j�J.E�8a����.�Ag�X��H4W=[R��������;��h+�a��l��A�aɅ��b-6)Lx7x'r(�iyr�*bP���	�	��vu�ip��g:� 2��C���~�n�e5�sEH����݂_���&wg9iF=�U-��m����6�D,���G�T��3=���="�4d
	H�� ��YH`��1���� �C^��Ā3����m�&;Ҹ�]�*�ʇ�R�	�t"�H��;�:���V��`�0�(��|����ͱY��&�|�"�I�T:��@�Q�̧Q���M[���騔��
 fѲ0�v�G=���O��C���V:�h�ZnY��<����$�P�R����󩘒#vk'�j�3���ѪѺ6Ҧ��A��ŋe����*j��B�������e�=�d i�P�s��L� +�Ԅr�� �.�c�f�@�|�x�z�8IST{��������5�Ή�~�)ڋ}nh}���B�W�;Z�N�����b�X��	F'�D[
N���
E������>�
}����,I�]o�?������p��|�({tm�h?sL����]�;e��Ȱ����*`�%;��6Ia�($	��	m9���%�	Mm�>'*2ҩF V��(Ŋ��0�X�d��AI7bH�c-�3�ɪZc�PP�W��t�]�<�6p�S�l��&)���;(���S K=0*������-0]Ow�@�{s&[&�Ж����W��x��̗�ߪ�C�'����J�#c���l�Sȴu��T4��(kq�}�i��$1O#,MbD����b1+����+r7�d6��S���c��&��=��,��{��.�ȏ�|�X[��M)�97�Ț`�2�O'���G��԰8~Y���vS
R ْp*t���%����K�~Yv�Vt��1�����y|��p(7��,�Z��z�ؑ��
�Pr�ы0
�V�ڍ"ԈP����.��ZCU�$�hl�ރ�z�\b��i��B���D�N��q��DL(e�����ف+�8�ӧ��e
ōNe_SC��ع�pE�I ����/=��1Ԏ7�fܶ�~�Z��������ֻ!�z<�����o.h�iα��i��ގ���[|��Ӵ�=$)S���an�y�2�:��4�xzR�3�>q��8fLkU֨�s%Ez{o	���ؙP���a)�䠐���I�_����@\L�۽����zr���#���UM�kd񁚂��ܘ/�"3+��@�	E�٠�*;>���a%�@?9�IH��1������@L��Ϩ:uc1�z= HHq".�R�i{��_L��p����6 ��2]�S�|����V����[R�k�9cf�iƿ�f&����?{2��0,��V��h�nv�'�כ.��'&w)г���#�pad�*:�pXe�y d�����(p�X/�\J"��)aRЀ�b�W��d[���`����}%\U���}�bB��ʚw�5U���=�#K����Æ����[j-���`�ۢ��maŗ�~�+mq���V�r5.͢a`���=-�|3�zxh�y�\��!���� e�):��N���PaǬ��W�dH!��m0���oD:ʍ��"�����a�y�U��A�A'�yP�����!�t�}A<�1cƦ���\��Z���!��{��1��i�_</[�{/xI�d�)���O 59+����$8�|n����d0�0օ�L�y��i ���x� Ci�R���}��p/����=�+~Y�4���5��;V��;�;�pw��G�n�������x0f�Wo�E�"��N�5�g5���L��SE:3gQ��a��mAfAha�i��jc�'a\�!�eW��	��9��tflg.KL��َj�~M bLhkI���ST��!����C��P��Je:N^曎����\�!s�eD����ٓ�: ۍ�Qo���S�wPZ4�DP�圵�H���*p�j�E΍��S�ޖCJ+0�RZ�PH ��E:��<�i���i�@�A�5h����!\���4���\*E�)O�[��s-\��M�ĳ��C֤�6+}@j.�1��Z���qȂh��^&�vX.K��/I���M/�4���GA�<4���N@(��j��}E������h�>>q�Q*�zg��\=2W�^�����r���
�[dr�Ho�=����A�7%��+}9������3����T�W�*�^1����KNd0����I+崄���D�Qn���ȥu���,�Y�,�����K��x���![}����j��N�?�ں�:O3�z��u���]4z5�#��/'��w���[O�U�z
��p !7Y�4���[j%!ZI�D�B3g���Hѳ�.L�f�nE8��R��H���^��%�)�C��m�߄}�&���j�����!��]�\�>���ڜ�����3" �A�4�C�w������4��:?_Ar=|;��tƕL�����8L��j&��OCXwKc��t�2v��Jޡܪ2�)��rb_+QYq���ɉ�^�7�Q�%�W�0�,��o�>*��8�'�i�o,Q�4$�����r�\2 R���2���27�D�K��*����t�-n��b��OH��/�C�G�� K 7����)��{>G�.,0�s�݈n��Ҝ���~KnV��)��A��ג�YiH5�rȉ2���OtF�G�X�"����� �X�7����-��v2��[�e�4<�n��#���k�8u�YW��k�4 ��#;�-�]�&m�utp��Hu�֛�j��AM��f8_��<F�m�2�;����-Ed�S����@�w��r�(���~d����}x__�D8�-߄�X���z��w���Lp����"d7V�b'ۇ"Y�a�KG�8�Q�Vy?�����T@��b�������OJInaϓJ)r(�¯�4��e
�<�W�[�q4_���fAM��� A�,2!vГ�l|�$��/�����Z~@-�*�K�Ş��m�s���c�g����Ї|�?�"]�Q���l���\�����EHECg4<�u��v�P�Q�����ȑh}��4E�_O�E���wh�� ?׀�`Y�.&DjKe�7="ɛ��Ú ���亩{|�wk�Pt�_�87m�u~g���E!�$gˬt�������;/\���X����5�aI������&�O�%����a�iݽ��V���U���dpmo3����u���2Vq�($�m�1�����m!tM�@��a-�!�$C?�r�.tÑ�U"}N5Qz5�g���@��G��4��l�? ��-]}�KJmW�9��n�[�Hk�>�B,�H$fTys��]C} ����]kws��K�8�FiS̡W���.��=]�`�Ŭ��Fp��xp�}v���-�����Z�'ߖ>8�%1��R��fXQưJDe%1��W��wu�#��m�ɐ����zkӦ��{@:٥H:�yLj��X.A��7n�+�f��ٳ��7�C�:���|��è�������W|��oD %*VD���]��ڣR2���ؕ]���&��&�!��Ze�5
��s�
ZH~LX.˭��t_� ��P���]����(S��d��f2��,��3�;�x��_�L^$��C�3!�^�Ύ���롖�n����/��<u�����Ks]��A�uT�42�M�Cb��G��#ލt��D��<�gx�����VY����"Hs6��r) �\~�1���0J�a��<4�I1T���
��G��$���f��}�_m�xz�5�s���u��l�PB��Ð�Ҭ��%����}8AZ�z�����|�|[�s��X���gڂР���8�������9S���'��c��x��z���X���U�^n|�u�HJ-�69?H	m�8���y�/j�	E��������7�{Y�B���W"�j�]��jS�r�E[į�<*i�%����7�ucڱ7bǣˣB�E���`�J5��"t$��j�;��D:�Q�b*ue�M����ֵ�h�Ą��l�2P\��2	_�hIw����ś����o�B1�	��Tr�V�u��A�|�)�X߂/T�5Y�ꐭ)OpC'0T���
c~`�E����C����䡈nA7X�8�Q%?�s4�[����e	��"_��	�
ټ^�i՗�;ǂj��<���i�jխ�z�XM�{���n�u��$��{��ɏȪ@���o�	��k��OSU�x�0+ȾL��l��+W��,�|
��0���z7t5����Opݹ��a{vݱv� loQs���;@$�{8�g&�c���:�>���� `�zz�$�%M�F���	�
�b�����,Ww��8�Y��4j���LN�۟M�*�\>3�9J���ғ��M�I/[(��,Ov&��e�x4	�R�1R(u���#PQƵ�
�EA�Q�5����Xڌ�A3ЯUF,_���0�@!��MM��O��Tw�&j�l�&I� dD|�L��|��b���Ř��R��k�CR��&z;Ȫ8
���56�������?�\)G`-k�����PB��L��x�8֤�P�aZ�b���� W�E�jom�m�A��h�X�}T�?�ۍ+�z�j�zdգ)�P��3N��'��E&�y -��$*���Ɖ"HF�?YQE&i�wo����4�^G��>(�9�G��� �	��o^�_���Ď�M��Dd�5�
��_-��W×zq��� �������ᛸ4mT޶ 0	06�T������dL_�^�Oi������V����r2�uF�!晜S�t� ~G�����	�ANN�%�$kܝ������������՚dᑖR0��I�<|��!�b��y��.IRꩯF5Vy�⼡c�뛁��y�o�;�l��&-�q�����e/CN��ӬK���nh�L�G(����I�ųM�'1/Bַd$.���1���_I�B�t��Lyν7N.
��?�^�a���������pKcY����
�_#����jUGĵ(UJB�4�v�˟f��� �O��ob�E�&�,6;�ǚ�I��<��|����!"G��Ob�]�m��A�L��i��9?Y��Ȧr�L�$,�xg���6�Lz	�Ai���vI���wa�����) �c�7��~���[���"�6��-�3^��"|���jZw�M�o�>��C���F2la�:�n��>�������ս=�?+Z�V"k¯o%���r�B��Kv�����ȰiV㕿t����] n3DDmu�{�2EZ�e����9��%���9y4����k4Q�:ɴ������@*E�����p2V3b��z��l����{�LQb@��{��'�^���%��ҧ}��>C4�y��������Z�	�_V>4����{n�������7L�kk\�
��8���$F�p�+ T�p��4�;6ab�-f��a#��t����b�@��m�4g��@��5�8�~Ï�K�	�k�j�Z��/oF���yͰ��"Y����~��ɛ󢯆p{�+�Ǌ�I� =lR���y΄��e���z�\b2 ��韞YR+�v��tF�_>�ɿ�+��`]�"K��*.P/yu/��3�
�CF\l�si�_�/���x'��}��#����/�@}$N	�nzK�LH[�X����fA�`���;E���O�1�{@$���>�+��S"�9x�hK��!v���A�}�=��\�su�������zD�Z[甇�X���5�i��7~^x3�P~���_��j.��aU�:�2���F��N�m��J�q�k�:���*l�Q��������IIq1Zt�C��s}�	��At�r S�7g�;�t�/s�'B������F0 �}QjG��|���G��y�j����%�c�����R&tQM�8�� y���d��)3ؼ�k�u77*c�H��.%$�]In�,�)�']E�%��qӭ ��ϴ�J�7��Q=��q�x��EPtغ�	M+;��ফQ�o�UX;���c-w�q����H���e$��Q����<g�vg@5�%pWN�v����͖�/Q��䝠�Y�.�?	��^l2���G�J��5C���f���{��MV��q<X����ڞ���KP���@�g[��W,�4�i��ӼiZ��(WX�۞����ǜ{�Zy��<D6�E/,�mn�Τ�]g���u�1�x��*���F��~��>�;�8�Y��	 3�ky8.��$�I�7;�z�,��f�J�L�f�� �)�ޑ
Gd��_&�;L^�K!��fq&���{�c�a����A� eq3��6�n.`	�}��0i��*��D���2/`x��2E�9�s�ra��|f|� ��&��u��\��,���ʫ<�ȗu��A݃�Oy�;���C��o�ff�7W�?$<�=��^�e��1{���crZ�X`���o��Z��3�xcd�3��.-�Q}�I�Fo���U�QN~�EH��I���U�B��~�9���G9�=d��%�ik�5��u@��
�6!�����d��P���B~�LH��]pn�?�	h*.-��,�9�ԡF�Ѻ%]���2�53��h\dV/�7,a���J\u����(�3Zf��4qԒk	(� 
�����l�sЄGv3Cs3w����89I}��ܬA8Y2l�#�d6�$�Y4Z�S&�;�4w�f�lH�Țe�]�!�v����S���i��NY�����sL�=_�Z}||�!��cڄ��VÃJ@��ҭ��_ɬ�גI�HX 郵�)��uF`4v�E�sMx"��W�A�����)�5c�di���ӡ��7���K��ŏU2�3ɡN���ˮ�T���V�z�!�b��닟%�D���I�O�������c�r=.uU1i^�Q�s�H���[�e�����>c��	aY�ʝ�	�T]�#�mS:o�x�ư�^�dY\P���G�b~하\�	�E�'~� �-u,Ϩ�eKn��ޒS�9�&����s�,p>"y��q}�9�f09�m�9e�޺7a��5��{1+A��V��^X�7�nV��3p �.�������VM�BթlG�/C�q���J���c��<��FbV$�RU���9GAa��V��5U18����	5s	r���:2E^_�M?z}���� �S)�*��4~I��<]��^����x#8����������}�:2�@@,�ߓ��3IG}�r4P�Q�f)
�3�>��T���9���F��] s(U�M�nX.�,Y�i�{&��Z/#��}	��Tc.��AX`�����ev���;u�A�2������Y)SqDź����O^7HafR
{�Q��|��LMY(-X�ι�����V�l#rV%
�[v��^w�gS��ܭ���#G񎗸vP�J,����z71]ΗK�&7��4�0�˜!�}R��pq���FoաU���#��&������#��Z6�6���Pe6Y{N��߆'� R3��V�pm���>�XR�<�\Y=BNҊ(�+�	�ʅ�����aE�K�3²�o�`A�y�YՉ�Is��.��,�I�u���_�Lޢ���٦9����Q1L����|��[F?��}��L�sf������_f�r�`�}�STC�jGUV�z�[fn���jd�.HO��+��ГY����H	��*<=Γq)s�֕lM2K�������5���Y5�(�ˇ'���:C�P�6�W={8d$ʧ�Kt�.���A*��*k#~�<tc2�����vj~<��k�CK���ʝ�Vuuİ��d]cBQ�FT�k��2����@}VZA�� �&� v���y��H�Ebco�& [|6G��k�:M�NB'����Z`$��L�jP|3"r�絅�A���T����r���J�[�#���*��u��Q'�"N�I}�{'�}�}xzVtǬ�����"����{BD]�~S��7|��ƥ�
"��H��Q���5/]�?���Ko�f+���-"7��`2L̩
�D�����G$3�E��!�XP�/�5�qo��T����ͷo�� 崳�*��KJ��Y>��-J۩��f���T�%��[�
�J#��w�����"��08[$�b�Y�?�G�s�ӔZq��ժw����Ix�zB�(��Ṛד�eR?��3��ㅺ�yFcO�����a�1�n�o�Om9��w���@�6B�Y�u��if� �ʞ�����Sw��Y���IkT����-@�S4�@���(P� �<�+��3��!�%,�������y�3Co���+����9v]Y�j�d�78����}�^���[�OE��{�.4
`>'�=�9���f�%�r��.(Q:��O.;&�|��a���"��P@lO�g�;�_~����m�݈��C���8�0��j�(��%[�IDj�Vٸ���Er�B_�H����Φ�݀��wǶbG;��QOΥn�ޫݞ���Z�h���`{��P{N��|��nsM2��w���8�Ȭж���m�`�g���Ä��bC���d�K�ܮx��c���;E��72��v�ߑ��ef/u/��� 3�����1{bJg��*y/T�+_]����_1�O�⡓ݐ�I��S�U�",��i�����*�ՠ���]��lZfϰ��_���Z.8)����_�a<���L
����͈@il&X����q�[ݤ�*x]�>l��
�c-G�6�1/�s�\�h}�hR�sZC�t��lz���.��ds�Q�5�ۖ<y��?���]t�p�"�4�#�\��\:h
������+`.��sz���C5��&�N4��T2��'09���#+�G&�qΕ�	yf�-�4+PR`N�(#�I�gN���a.l�)��>��XMJe<�?>q�r^/dx"���1�M�I�jY��8�����v0��P�cS���S��H���=֮��Z-�a�����.�1o����$D�	t[�H}t���ϑ�1b~VT��-2\;��#��WoPL]���Kh�Mh&�H˛Nsp(���h#҂� �z���7�)C��nq�����jާsS��h�l5Nʾ�2\tv�aֽ��-���&��v�� �U�{��"�![؜�ުD��$n]|�ݻ{������}gkǪ��j��+]5��pz�P�},o����6k_JF�%���1�[���4؆6��fT��Na��|�����~���p$��ތj�,[\��F��yP�H�r�T�(�j`�66�s�=?#��_2��*ho�5��.�C���&�3Urܩ�����I}�J[��q5�?��xB����]B���
�Ip�S��(K�<�ZY�[i��ɬ�J˥x?�� �	t<����d+�N3iϲ�_�}D}b�����F�`"�Rp�Y�`��*��0�#{n>���w�c��E-�=��3�sqXS�b-�<y49 b�I��'㔅/��<��t�����d_"�+�'��|3s�X��mq|�'-Z�bJ)Qv��m�V�����S�W��yߩu��tS'��r�}m����Ⱦ:A��P�`��l�P��\�"&�PM
/�c�Yt���&��nO�MԬ��^<Ŷ�*{��@�]��� �Ў����R��+@ ��K��<gj����br}�R��t_�A6=��7����3�Zx�-���ρ<3z�G�FkY���eEԆ-�d-Ů�$ϳ^�����]��ZD�������:"/C�a�S��`��UZ�r�|aͦsl���������JVkx�4ŦoƜ!a�S):I%�����5	4�&���u��Dqv�j��.�G}��aeb^��)F���%X�hmOې.6]5�������r9٘��x�+�/��$�l�:Rn[�=-��xet�B�C�0D�Y�=k4���=P~hG�X�&�D�4��J���̻?���]H�@>2<#�������i�j�y�>KnF�e��a�
#�q�C|��] Iv�+��d4��f�q,@����t�=�9��Xd�������ڹ���G*/�@�T2�;dt
1�1�a6�l��*���%U��+ԥ�\2-ٓ�T��=����Ä��S��MN�.
�����9�Y��h�s���<�?���V�2�U%d?�:s��$�#!��%	&�:P����w�_��+�>[ߵ�_�'|՝fߌ�}�9������s��zhғ���6��_���"�z�E��2�Җ!i�y�yJ,�ÑoʈJ��QӮ
\41����Ӄ��Ȭ�
7����8�m���-��ͽ�T��h�[�X�q�A�ԙaxa2�W�&O9|���pAU����'䝰�1y�!��:�
�3��%zlEl	�!��v�?Hܺ���&n��a{W>�Q/q�_���%9�=���:֥s�@��f�I2�����[�-�D�C{h�7����0��j�qւ6"� K��"A�G| ���'��_�8;eB1�9�PdYq�4C��+��>e�3B!8i#������ E��Y�	�	G�+^4�V�Dh�e�7߼@�#Q��]H$.����:���?!�����ץ2�s락�h��yZ�L���s�Ѧ�d�A]$ռ�[C�D�s`k��Ng*��A�J�8�b�ޙ5MȘ�O��<02I-�_�|�zc`�ȸ:x)r��P.RjŊ���,�4,�sK �~�mY��I:&]��q���I/��삹0�����ۼ*��{3GO������[�Ħ)�˹{��/�����x�?`W~.b�'ωs���ٌ���0�P��a�Ǐwu%5;�@V<�<�޾�*V�e �{}OӜ�	(��
q���=l;���ErR�H�ܥx4��2��1��0U�߷3�k�kiǻ�����}t$FNA�ʘ[.��|kЇ��&"�{���_�,��k�A���o����Am�A ���#Pb.�
���I

7݃�e.�%�8�1�2
��#Z�ХƁ��6�GdiT3�	9)!��:��de<�Cl��)�7��w`��I�L�)FAsi�,_����1���k2��B�L�];%�����,2΀���U�Ȅ��H�g����j���<�����\!���$�h�-䐛#��<?�!R�i����
e�[	�y�����v�{M_u��EJ잛��p�.4�is��p��rX�DO�'kD+?k�]�ς&�� ����>$0��Cu�EK= ��������e	f�b���zK�(�[p-�[�Ѷ���&��;
��^�1Hif�CV�����e�h�[���$�!iB��O@:b��`s�� r�q������K����映�-ά�U�/��M����3-��r��/�2�8�>#���{ГqƁ��K���uG�3i�6#�j��	�,Л�S�7�K�w�/S�����Kx�x���+�!Z�VMx��n@MP_���9��2��ֺ:��;�:�,\E�SmE��1=D������`�Ѡt�?�fdtF��0`��>�Ը��sl}L��T�]QR:xH��٫���{��8��]%0��Z�$Ȍ�v�^\�}���O7O��mc�=�@��o�iu�U	D@��X͍W�at �����Շ�iL.�W�(�����T#u{� Ŀá�u��>.x߾�R|e�`���`�=˸�����5��W��18��.BW9���7����*�����%�t�O�Rb�3<$��A�#cD�'��3�7�A���
�硂h$��m��x��EjJ&�n�i�Y������y�5pw�Q+�"u��hH�+�LFm��}d��Z͎%���:���ĐR��bA�k� ��yQ8R<(eLA��6g��6���עP���E0g*E_2�^8
�Ļ�!)�3�v4\I��P�l��V5u�����&HV���t�@!v��ǉ7�<S;��A�x�n <�J�S�؞H��h ���[e�w�Ԥ��� �0��H�aCJ�M��~h{�~/�e+�f�>Dٮ\��c�|��7�.�%G��+9����wڠ`�X�Ɣ_�%��E ��S��(4�:����e�%Jq���͠����;ӣ���V�J�-Q�H�Y�ܝAT�������B*H�>����9�X��?�<����
Q�̐ƞf(��eB%���n{b�-��Zy��a�q���)"0���A��

�����WY�7��@!^��ڴ������ Y�q�]7�5�d���G��c�󴍏�&ł8�߹8�; �Vd�f��'M�G#R/���v-lY)�G��
У{�y��Q�L1�)BK�5�L/'������)�����e���
G����<�z9���J,���J�{�b�C�B������f@0�Okx��H�Ey����2�o|�C�f�vR��԰����ҕ���E���A��SI]A��]���OY����X��J���4�(eB:�%%0P�����5����~��³��II���ᰖQ~�9FF�h˺F����n�kn�q�F�u�Z�MGp��͠+wd�G江6���VOt���22�fI���a��?N@���AG�X��:s���o�9/t� р�����`��!�Ձ��N���#� ��ﶟK�aG�{���f�u������E{�|r�>,�by���S2��`F�FQNZ&�K��#3I*�XH�T'>O#,�}[�= #T�>�#U�g�J��*(���|3�>_[)8l���V���3�Ҿ�&ospp�$4��i_��f|w�o,����l�\�x�;~-GI�;���FT��h��6���ly5=�	��E@t^��O�7�b�(d��M�T}����d�vW=0S�}����v��E%~�������Ĝ�	�q7��.T?jL g���x�x����{�����q�}n���LL1"��9��=eҾ��MJ_VRe���"�I�����K&`�I���e����Ҕ�k{�-�N@�'�D+s��ٶ��$��m��Y�%B�`���C=���9�������_Z�|f�l�o`R6��;6#pDn�w�/cI7U��EQ�C���U�2O���v�Q�0���l���6�j�d�vm�Ը�,rո˜��2J��e���t MoV�І�O�����~fR:�����/
�;4�Lۀ1g��f���"5���D�հϗ	4w�4���4Zi�}ǣ�Q���.� R�n|�
nV���1&e�`	Ko)��V-���˩7C��-Y�\�	�"�/E�,�6'GA15Ah[����\��E�1k���A)��֩_ x��7�Ǚ����=��ZeYh�o�_Gb)�ϳ�s��*��φdȒT~|��	�^`:l�Uw9(}v�.N�+s���'�=\PG԰$ܿm���aQwג��i�`<:5�2��D)�����ڟv��:���!;+ä~7%�~�����H9ȳ99����d��,���J�iA�	�Z@���[�O�ay����)�"�[n粦f�s�=�����>o�@Y6^�ϩ=���J���G���mɊZ��#��%���)K����#�-����\�_hj�ԭv� �:G�#�����D��l������������E}ىG�������w�QB@����)�
7K���G����0�3mO� ���JWH��<2��g�,�Is*O��bcZq⣒u0�gs���Q�7�_cf/�x�W�e�־���\�Z��0d����Q(����p��Q)sn���;���y�!ߟ�k?x�����(��r��)�6CP��x|[�����\���9�7��� �O��ܤ�����!��gf`�c��5��E5��8ӊɃ�eg��������%F��8X��^p��9~�B�>�f��,%�~I,1��"�K�����iS����(� P�w�ȍ�7�P���a�ݻ�J��o�
r���������Th�t�HQ�9"x�8΀O�{����A�f�Lkt''�<��+1��Z!��('D�wku	���4-���'Ī.�r�-ps�{Z)���.H0��_�.�c;R��������5��(���c�뉳'}�55A+8���-�,���d	t�j�YUC����C�F�!s�xH� ؅�K'*��̥!_.���7~�ahq�*}�Dĭ�g/I+P(��2؂��촪�̑(�����P�d�^�t��W�:ɠ��o�?7�a�W�C�������"!�����S��~P �>�𦾧�xW��fդ
��x���b
D�C�@?�JeV���d��@M�fY��
�*
he��"��ބ;�������o*Y\�$�$�3������08�#M�l�%��#������cI�E��H/�a��g}*{� z�����}�HT���"/2�g�m�>ۖ��3+��!�?n�;�0�d D��<��hy�X3�pS�)� �.�"�T�B4�Z��q��@�v\r���:���2�Xz�A��̃�܃֖7����蒱#M�HX�
����9dPBUoQ;�o{�+�%jh1������!�˒��w�
:5�1:�dS��禯�B�2=G�+,qB4@��֭�7o�܅��Hr�\DS�� ��{3�)��Gx�.�tN���>MJ�Y��1^R�w_��^n���S�Gl�C��Qy��s���H<�|8�����>?d�iٵ���x����� ��31�y�者����gm��T,���1�����]8���ss�Su�_�f����鄪]qh�@n�@`�m�,n������M�u��C��{i���dx�W%)�i�[":CHq�п��Z(Tavg2�hmև
����͍k��� KGꋃ?�v��~�x�1n4�W�`����Ŭ���m
7��y{h�V+�+q�VX �;�x��8T��%�U�0�@2{��ͱ��Qg@l!H�R�'�5�X
rbg��r�f~^�c�0�hh�G8b&��ۘ��'��*?"�g=�
�ueLd�s�u�m�F�xH�U�n�3kt�9�I�xǷ�rM�;�ZNJ�::}5�u_|w)8�a��B=Y������C3 c!͔�1M�q�~UX��%Z9Gk����`�b�-�SLYe��~���ְb>Snu*xgP]�7�lƁӢ�\��}tG� �4y{"�A���u���w�#��w�:d���;�o�_�����&�D.Ed��y�v�(�ow4[�e+@n�K:TbŃ2GK��-���{��ܮ�+Ic�I"~L��	���)8��}�S�V\Q[Y�{'�K�
Bd��N�� ?^K�7ТH��H���`�q�s"��X�'��g�+5��Zrb����p�����q���f<uF�s;��lf�ŵ�lj�T�}��+��+�М)/���(*.�|	]~ή�D���,4�!�2t�҈ܝ���NX�B����ԉ�ǧ!���E`ћ��y�&a��}��K���d^oZ�p��du�<b���\ �Y��9ޚ�������)�\˘`<ؙ�� ����V���79���I�;���i`�vzcO2��w3ey]��J%�]UZjيb	kF��*�}��]=�ʹ�(�%��0R|s·7�{u�NI�+E�ULFl����/z�
̖�ng���.��W,�O�l�ԇ�Z�M�ӵ��,�2�4\O��qeLM�
�prN� �KN/.��|�����}L�x2�|�N���������s��1^eƫ1�/Daт�|�x�z`�9�_� � 4���kK��+er����v�5�m�dk���)d��G�h7�	�����^Tór�R8��9�Z\Q�i)����F�Hq������Y�೸��:���trgO��!�S6�v�uSTX#Ϸ��T����B]�5Q
*��C0���G9����7��'ʵ�4r�i�>��k��l|��0�Q�w:Z!*�*k"
za�L�dT|%�v~
]�h���.�YVQ���J!Ky��?(A[¢�'缰?��&���[G~YO�"^�K
��ӕ�%��㐮n&c��C�uֻ�JT?�w䐐�����Q���txZF��`ŗ�� v}�4�˝4�] �i׳6�Q���8;Y%�1�PR״=	�E~Q��2��;l�/�~�*mJޣ>6��u��_�f�1*�
�����Y|---���o.�
�o���A�k�c7�)��֚����E:�X��W�r�4~,:[�8_]K�<���"�řo�9e���x`����^K������c�Wʄ���s
��]�� ������ч`6f�z���\����=���VyY��p���I�v�=Mt�[V)PA����b��={ϩ�T%��^�0�V)ng�B����Vx�w;������#T0uD7�$���{z��*��|�hZ�^S̃	 4�L<,[��n:ʭ�V}�kv*L�d<;�}�.㜓�)߅E\Ju��6eN�E�}L�� � �+�P�R�z�f ���y߁��ì��:��A���v��C��	VA��{�L�����r��x�0*�w9�=�6��F.3k$��Ȉ���G��+��mI��t."<��;uMD�Amh�Cͧcӓ&)Y�(I�}_�z��Pk`�6��/��[)q�X2agO���Dޗ֯b�k�n�>׽��`�8ڱt�zR*,��*>
\JF����"w\�k6��x�H�Py�8۸V[TjR��T��"���k��&*-�jt�Z��W��VHX�FH^�_���-�z0��,�����U��%�V@(0Bax���2����>x���?�S�g-�@eB��F�M#�\� mr�5%�X�U��,a�n�1$ҩ\8cՇ1ά��(s�(,k:wR�W����Rh��P��`�DK�I�q9�>g��B}�`R���t`.�u�<?	E0���׼ĺb ���P�������Ʃ#ः�m<Z���o[�T�8��ygj4�fv���_D*��|u1� ]��p����ae�9��ɛo�Y��q�m�=���ni�$ʵUt���Bb�Z�襣��Ǎ����-��5����'�>YP�i�l��أ^v1��ѓ�SbZI�-�>�hY�y?�.���j~��ѐ-����������Ce7�6�>�4 ��oHP�����N=�6��mF]�M�a��X��`}�ީ�	0����4id@�������KVx����z�D�]��Ա��)�s* j��>���;�%� }��lOED
|%����5�i#�%�N�	|��PLع��V+APb$Յ�L���2�Q�����TE�QTWSS��\zq�ѹ���B�x���9WCO86��&��p�ֲʹOB��S�3h�?�ρ�KjH�L����d)K�K�5��nn�Q띵m�,!�ZYi�.v�#C��+?�6�`�+㩿؈��a��bk[r܋IX�s&>m����hHHUɮ(f��s��(�� ���	�<&#�
��������a`��gO{"{����j���m_���]!*���B#�`#C}G宄��l��Q�I�h��s�ܚ�l������6�O-�h�qߗa�q,�ġ�
���.C��*��H�����$�Tmw���4�@��a�# �As��$N�$e�Zk�rP��Q���/[���M4k�s�9�
[d�J�Ȧ�(Z���&��iA�Aj�؂�Y]�y���S�t�h:4k9�������X,�5�_sT��s�k��_#Z3.��ϵBDQߊ��`j�zx�tɋWjJ�ڎ�%�h��|�Ո�-���2���Ұ#��(�����6aX�bι3� �$��G�3�pQV\x�7m�gz��k+������hgIڊr���J����zXFg�V�%���N�n���$�;��m2.m��U/����E��˗5�nm�V�����R;=>����J��}�B>]����;vJ޼=���E:����t�ɴ�����)�Σ�{�F�X'G;2� �+�I���ʃ5G>s���6�/��#��wY��&=�I�"�=��'*��,t�\Y�hՎ�`Y<��Kq������=��>��L��4��xT��Z�h牿[$��$.4,�%~��q�_t���d�T�&�k�Y@Pr���%k�O	����3��J��r���cp��23����/m�� bQ��K�	���խ�K�8{�w���~d���*hq�	 ��������6�A��VC�č0B3F�o�~\nNJQ���'5����zS�[�2�)	��/�uS�>�F�	��r~o�6�]M��͟�[���;�s,6�<�>�����]��������� A׻O��Z�0�u� �����ԘǴ��i�k�n�o�e΢�uܒ;�0�d}p�
�'T:�'�*��#$���ۤۥ@7�)���p��.���d=�?����),�������d�~l%H�MI�w
���Jg�p�ϓ�[׷�X>�hQ�Ӑ w��O�b �)�=yL�e>�̑��c+��&�H[Y ܿ6�������&���L�O6�x9'Mi)�l5�X�VD�[)��K��$��xtv�{�M)=��Ri��ե�#��f:j�n����`/$Q�S�>���Lm������FT�eA�n��͍.H���:{���mma>+��8�o�?����4~B���WLG��	�ޔ
9����)��I/���qWF�?A�F`s��4!e^���7ώ�Q�Y̷ؑ��J�T�r1u�$��A�<�"L9��d{�Sˍ�}�i��=\���EEZ�(#�^�7(�;�ѫK�/�H�ȃ*�Y��?�HSz�W���g�?wՑ��u͏�b���C-]4���2{b6�`@E福;�_�:$��FU��#� �5o�E���?=!1��LmJ�aw$��-2��Od
���G=��X`R�W�>=(�UfU�
�Ќ3��婀A��N���zX����������m��X�j>ьEm&�AL�P8$`�/��l�,���u������ZQE�k�hȾ�s����H*iT@�l�$$���:��pɈ�2��U=,�΢�6甲����G���T*�L��N��,Y)�\���Q��N� b᭠�ޏ��q�1��7p�r�òߐ�	j8?Xxǝ�*�~>D�������~�:`� .O�cS��O�v��L���a����%������y9B�.���oo{t4K;�uTp��ȠN'\�Z��7,�,��7��Ϸ	K�iw�DW�b�w�?x2&>nc��N�Z�J��4�Yza&'����%:)�w�K�N��Na�Y�%�����L�]���{X��hZOH���F{�X)����hIYx]%�t�� �˿�1�@�L�o{Q�<���c#�P��#��T��������y~�F�A�݂�lq�dR]í���*�jB޳&���B�ަ��7�zE�'0;av����+{�?�!
���6�����5ՐŜO�Uf���dl2�?,�� �)���tSG����~~�k)[��y0��Q��]r<aY�7�����@�4I�����D�ܕ�P�f���y|�k��tJM;���ۥ8�8�E�6r҅y8h�<�-<���U����4!�{��i�=�-f��H,���ٰ�1�0:%�ET)K�"m\�
�#ԃ��NW�#�����n����"2\�3�ݸ��y㑛_j*@yG�@����^���c�M�����������B}E�z(W�s���5�|B�Z_m��ʶ(n5 �"���9���&�v.�I
�0�n@�g5����, ��A����6�=)��r<b�@�%�l�g���|�.|��8���4�k����0�T�ħ���C=�����3�qP$>��c'|{�<��K�΢)}_N|N]D �*��������r��C�љ`.�Tz���ɚ{�lP��f����tzb�x
>C�Y
�w�܎,���O�H*8֞g�T1e��8Ѕ��9�	dg�����`�:�B���"�zg�,x��j���5���l�g�7f��x�f��Eѩ@�����E�^�ܷA!�v>���o�7����^�P�2��V��:�����V3
�vp-��WG��L�,b_���/���*`�}�c(��� sr�]9U���_xċ���`���p����G9}�24�a�BQY$b��Y2ڝʧɛ�ǒ�CT�Ħ�(,����=���5�U�� ����F��FY�c7,Y��zc�x����Sr�)U@����i��c~�=:/�1A��ӏ�v9��)�_ ��DZ�e6�vRCن8'xg�+�2��:�hyѳ�C-X����ʇnTj�4��XF���4x���^B���!1��Qo���)��0_Ϯ���"�� �/�N����C��Z��`x/�ݶ3y�!�ɕNapR���?^����3f�n㡕,j*�6�*c���ڔ���V8	��Ia��WD0 ����Q4B�$u~"P{`|8�K�2���/�w3������gm�I2��%{�ț�c��`�$��N!v��Ӈ�6Ċ5���	�o��P���U���6g�p����;�\.<��:c*(�s�Q|�zQp������J�=UB<Sʽ��z�
�������[��� Eg�^�n[i��NW��ɗ\^ �o;�1�+��qv!�T�Y�A�A�}G}1FG�A9z�C��t��v㧺i���༞�rkFSF90ig���x�Gdf��yhB�O�N|��~$��48 6�H��Ĉ�] ��M���冲�ʳEQȣ�a�(/��_mNwEª5d��|&)B
��r)y�.\�S��C\�*٣��^(Q�9��8Dr��������Pa哠/�_lP��lWÐ��kiI=#J���򵤄-�����q5uDr�N��(�P����:,~���X9�Bu�s�)D��׺Z�C9~,oM����M>B�����ܺ�������vX�c�%�Y�q��>i�`��n��,?|g��.�4�b#}y��˸��cK���1�w���$Ez�$�<��,����&Y��yJ��T��Or�ԞV�bdr�B}�'�}�H��R$;Ɩ����m/�R�î5	��4���0.��	�	WM ̤�N@�VAwh��אR�r�=�t � �h _��<�4��~i��ZQd�'�UR*�#7�i��$識-Po\��(i��`��1pBҲ��e�C��l��D�8Lɶ;�c�{nF0j;m�(# �P�>��MᏢ7Q������O�u����#����=�I�0�`ZѶ�l@<�҅�'���E��ɲ��D����s�3h&#?���F{j�+���İoMeϯ�֢ZW��S���kD�0j7�$�z �0��k���;�S����ǡ��s|�L��">|?�v�m��w�T�)���ds{N�g�+�4|�������$*U�h�O�����r�/��q}"m��J��y�Pݢ���
���)6:��ѮP�2ah�h˯�}a۪	!>A6¡)�>l�b:JA8Ϊz�H0�"V9�j:��]׈����g�d���gڣU?[��f�98��$�~���zI#e��G�Hx��E׆6L���S*ړ���e�_����g��T6�*��d%���(3C
n1���X
 >�X|�)��EA"��N��X�fɾ�E#xS�i{1��0��M��pG;F2_(��/-�=k�3��[w����m&w%�;��&�f5���k�@�D���/�T�)��Cn�y�~���R��]��#Xଦ�
��p������+S�p�sK6�3�^M�ݽl=�z���ٸn�:��XNl'�W3��D��lM`�<��0ÊŹo�6Sp����=U3y:�� eR!�Oc"h��Ls +l��Wq[T�,11��w��Ի���S�u*J�o,�a�t׬ܥ�l`k���܏g�4K�������>l�<��@�N�k�,�9Z�|~oTi��/���8'a��e��9ކ�Gxf���j��$�ä�y<��3�K�����] �DL�|��3���Xb���bB,G�'�jM-MU���X������v��	��C~����~�wN��l�`�:�x�-#��]Ah��n~(�z�l�W
���'�OB[*x�T$0)�X$�}.�x����`�t�â�����%>�'n6����a"���o�+���/�������?q6�h2'y�õ��OD�I�T��6��hg���l�f9��`�#횖#�@�+���M�c��j�d��g�@�/S$<���ӄR5���<�T���3�x�]u�iR����%�Zy	���wJ��7�{�ٗ]yH��a�f���h�'z1��|�"|E�#��{���+�9����f��=J,��K�C��'\��池&��n�����$�
�L�&w�8I��o���VY��}F7m=�f*Z(X����]���f����>�ms��z�%4����?�5�����K�z�ѕ���O�׉��X��$$���SU��4v�Z�(�@^ǛD��E�_��
jg4�R�'b�I?�1�#��?�GE?"LU.z�t��Z>��N)�1Ry�vҤ��P=T�9�ry�-�E�>;u�����0�֥-��%�v*65�L���Ϊ��g�@��rafJ��jw/����4g�t�{�'i(�$�N�#MU&W��0D�� �t���{�%���7�wjn]tA�b��`�%@`g���%P�-F��AW��/T����	Ъy�_�M|=@YO^n`_&1�`u�f�O���A�ة(�M��v=;V?��s܈]���(ڻ3E�vyj��vغ���΂����Q���{���:j��lھ�$a�2�Ǚ�a�l�A3m& ���g7S�߯ͩ�	�7��uL '!���z�0Ӛ��"^�M϶mb�ł���O���F8m��Ш?%�RC8bP@T2�F�>f�¨U��b���o �3��!�z�r� �pSI�!s"@V+��wim諌A2�m��s��{ o*� �e��������B�	� �Od�����}X�O����e�Yz���t���q�l;)���]Ff�^Z1�g0u����P��[�Iq~��]�K �����y��7� � lү�e�_�ـǒs^����Q�\1P�ZOzF�S��/&d`;��K��`)�Fꑫ�Ue���';Ї�I��ؔ�}t�p,�[�z�B(�ȅ��QJ��h\�r+7K!+lt����� ��8��(�:Jy���z'�����f��ݯc���%�����y�d�V�b��}`��cѵb�T6r+�]�£��R�9�h�*��� z�I��7�^l���1��9����4�.
�X�5��C ����0��ShR삽�bK�r�������$JV�O<dG����s��0*��r�+��qmh��f
��6;�ޗ,$��Z[�!�!׀z��1Ǵ ߧ�L���A�	�����t���R�sV�v�Zal��Q�
�uW��<c��u��ܚt"F��X� �pߪ� ����(��(����b~�Z")_oQ�+� *�ּ[۷�yQ� n����,iN���wl���P�D�?E�RBs��>R%q�.���������l��?��M��u�˼�?*�I�t��?o�H��<��c��ۈ�I�aZ4�Q'�����l\l���r�hm�H_Q�p^}��=O�Q���y�셩�%�pg�>UP5/��|���~��H-�QX.u����¦��L���x�V��r1�j^`�/vޝ��"Җe�d9��J7NiP��?oGF!���}���Ny^2=Z3�)x��Pg/�喆���ѷ�������!�I�8���H	��2B3+�`f;/&��G>�!����P/�$��#��
,S��B�-=�D�Mf�l�B�����i��B��6�@wnvQE�Y��X�I�&�-��������FG��LE`s Zk�K`���b 
ͷ�]ְyK�d��n��%<V��~-i?��H� 9t5:�(�4U��{�5��̿����L&{ ��n0;�Q�
��ծ ��#(/��(R-d���z��9��+��wm�40�#8�˪��Dɰ����D;`�t�Qt�c�?�hW��Ȣ�y!4���O��3���*�n�Y;ɾ�&(�i#*w�9yVQ®Ѷ�-�).�RQ�n�Ru��LU-�W����w�R9C�e�x���Y�N�,�	K�`�V>ܯ�%9.�!��R�/�ғ
bjC�W��ؘ����~'���^�G��c�V�DڃI'��|��>���8��A�[�?$A�w3w�!B�C�7t��f�/MB��w���*4ui����)�#e��<��KK�d�uR0��M;Q������'��$/�l���^\�)
�V�W�żÃ����2�vu�����x8� w��Y%��l��ޓi�4g=� ���j(�,��\�"V(�n0ߧqurۖ\�vE���=��w�d�����P�Z�R�*>��N���\�;�7�2;���g�
�IM���yH `L��Ӄ�W��M��b��è�YR���zF�>B�oh�c�$�8��@��A�E�*����u��`j��Կ�m�^�ZLjE.#+�-X���0�H���7����mڋA�0MNV~���ȳ]��qg�Hbm�R�h%�Yk19����c/ӏ#���o]�0Stf9,x��Q���2ޝ_tZ���}�~|���	 ��B�?@b��W��Vx�X���J	[G���rMv�ȑ���r���ʹ�<��k����lG"��w�_�<����ɿw�tk�E��8
���˾蛇V� ��y�a���@�$���WÃ&B����ߒ�NT�W֧1�H������?M��+�GRZ����Pm�Hj9�&}yyȾ�"��w��
�t��tjk�7׷=;�0��t�OX �m�߻�/�uF�����֭h��W��W��s5�?|e�?�S�x���OΫJ��T+Z%F�˩.�2���JU����)R����ʥ��x�r�wQ<6Y�[�3��Y�����Lիʻv4c�)|�3Q�7@��9	���C��T����5��#���D��~�"&�7�h��=�>:k�nᑐ��o&j)�y_��j �\�7'tm��h�����ʥ͑�E�����'jv�ť.�\�o��#���=}��Y4X�/u-A$�ns����HQ/A[Ǉ@ϳ������P���R�z{Gb�NlMF��&��5^�T��K�'��L8�x�-e6F{�{�e��)G����=�b��ȼi!J`v��������M؉���V�����􎺲��Q�$�t\��9dʋ{\It�m�aO�Q�f�+hŮ3��� ݵ�$з����ru7��0��IUcJ�� q�v����_���-��m}��,c4�d8�'��-��.�V�� jG
)>G@e�|j�X�McX;Z'��x�N���Z�ӈڢ~����@vx@�=����%[��0�Ҝ�tɖKy�@������U~-��;uZ��]ĳ�E�kd�+� O�mK���ܠ[?�D��3x���H����&�7��3�=�\�{��cE:�
�rIqt�m��yJI��#�d�6�"1GJ:"����I����W���	���'E�H34���&f<�d�Ɂ�:�47��W��-���T�i�S�Dw�K~��i��;�X�y�������|!��݃L|� ^�1 �'W��A[u��չ�h��K> �B�@i�5]o�晊�6>��S��8N��G+���eq������~�y�6��ɏ݃���3���S��H�7	�&��~�[C�O?t�����p�ǾG`��!��+c�S{��>��X��![��|F�� ��*;��S]A��z �"� ��Lz4(
��q��n�u'	0X>���%'�W͡�nkȩ9՝@�kJ�SSZ�~��T��	�S�wS���<E��	]jC�-��'��(��=b���>���P{utr����Sݵ��8�ϐ��@��I ـT�5J�:})�	���.�.��L�0=�"��/`/�Ѧ,3��ZD���t�D�nI������vM��t`�M�(m&��B7�7�j�4��� :��\6�R�%qe��J`���|��Z7y���I|iS��kO�� ��S���0�<�a�n�f Z��c�&KW�L8pۊ�=1�
(�,���E�a�.��hv����꣨��w�u�}K[�����M�O�t�i��b7�~� Z�yu����ī��4p�d�XE!-cn�H���,���(+��"G�V��L_���SC���W�̹|��d�ŀO
$Y_��w+ �݉daҖ�iԴ��7�P��/�IE"�c���L�v�Oh8h�:p�H�2��
m5��0s�x�豿�y߈	��U��/��7%�(d�\�|&��|\��ɹ�<�g�e@YZ.�>�?c��hpN�B�x�A��W�P�U|5cPІ��W3p�h_�϶m��5W
V�1e쟖#�������dp��8K��T#��p�
k0�vk#����.��tL���m0�3ғw�B��v;�$���.�d�x�]��M➘Oxe��u��p֘&,V>�P�^^�j�*���j�f���݅�jNɣ�h7�4�;�D��.J�5r�l
V�~YГ���	����t[3�tE�C.��3�}�]dV�J]ѣc��R�P!��D?������SϠbkթY��؞�4zDΉ���W��� ���� )�ʹf߯9�'�B��ׂ�f�� :����m��V�0-.[	'��Is�=>1������K:7���4��u�R�2{-�kf2�d2UJ�Y�u��J` �;��r����V�z�ԣ`��0����ʮ#�뎷���,���[	5�T�h���\�]�pU�kΈ����Pn]�ץ��<��f.u�t��zo��
&�� �9�9];��I��	Q���+��m"HJ��M�L���G�#��A�n�������4�q� `�c'�ʜ�obY��������z��(��ϕ��!�ocI�֬��i S)��Δ�*�(���?��-��W�,CY�R/�2>�&�-��Z��b}������"�1�@���Z��������f�U�a�MFT��Ǝ���Y���4�^Jl�Z��a'eL�h�6����U�[Pq[a��e�Z�B��s|£s<s�àXoG��A����a)RO˫<�ܛ�� �fD��ٜ̍A�iLc�6e�t����i��t�A$��:Y�����A��"��eL/??*v�!'ގ�z�JI�X����YV�f���2s�8�Lݻ"34�F�O.�k���P}���+�3��mn�4�4��d�Ձ�酄s���.}�G���*'v�ك�bY�`D机����0���U���>={$|i�qt]s�<2w��Ѿ��1u��;EB���r�@��ߍ4 B@��6���*�`	;���nt�ϰ���� �q�?��{��!�7���͘yJ��a�W�԰c����$����0�)�*yؾ+7xl���Ehu;kX�<KT8����/4�@��� +�Y�g�t�zh�GwݭPt�3:���*�$g@/���c�9�P��4Y��i�N-�i�Z2,!5��G?��z�g=F@6��<>ѣBt�����[o��!��ʡ��Vg-�ə+��b�TUsL=#�������N[�J1Ʃ~ �a���mBG���Y*�p�XS-��}4`$D�Q쬳�O�m~� ��2w�v���$�+�o�h�x��kk�Sz�8Y�;���A՘�b˯ˑ��0#rAG�������Nղ�綧�{����|��'��y�z �XC��S�,#���"��f�
��t;
�/I*$�v�78�6���D�}��\ :E~�H���+K���)@sp��Q�����}��e��A=%V�1i��ݠ����w�z�O��m�x���'-�x�hк\d��������H;z� �'��F��|`Ђ*:��b�.�����?*�hG�嗗#�&� I�d|����C�@�Dp�{{�9�zJ�PA"\T��ס1��ҌβJ<�繬�=/�R��Am�����K<�&	<��Q���H[���>�3����┐��WUĦ'~r�l�-ߑ����Pn_8�tX��O�3U�y�	1���1Ă[��=v=Il��y"aM�)xG�Ǆ��J�+�W��%�j���C�r�SBW�3I�(��㻭�������z�O���_�����*����p�ʊ��W��P��n6� �Jޫ�A0#��1���3*�"Y�΅�2ה� 4�z"4��	P���z�$�[����d۫,Mw�+[�ɬ7M-=LjٸB�cКY�&4:�d�ؔ�[�qq�ڗ!�Gc������s�~_%-s|#ؕ��ýha.��o$rd� �~���}"�5ڳ�������PA�G�	3
�`��!՘��R�P�1T�S���)A(j����؛`��2U�6"/'bc��m.��+Q�iF�a��ɢG#��+�o`?w� �QP*Y�܁�,fp�ھ��{������ݧ1��e��VXj,���F_M��_��IKJ�Q؟��J^!�#n�S�g.�^m�F��(��?��!����*h#-I2o:I���ɢ��PJ�7�v-Ju��V:b˷mޞ��8��~��v9����N�s��~�����s�������+�����cIo  A��ް�8_[���G�F�����*1ӂ&Ĕ' eP��&�"ʟ���c6�W��i�`���,ԑl��*�\�v �x�u�[��Z�!�� 3*>��/�i(��j�����ۛY5\�`3X$%����L��4WL�ȁ�Ǯ)�crb�ߐ�\)�LV��CK�����	1Q��x?����4��vU��!����X��_!���I��'�_J���̍s����A[5O�����m7�e�9fH�n�ҲS�(4���n(�S<4y��w
������]̊�hAb�+3�*@O<�D�B�0�2��GD�3�����3�V.V��\{h(�X�O�BaR'����A���k�ɜ\�%�阐�~��nBm<K������P�cFCs���7���}���[0]-�9�ʈ*X�vZdȿ+򹽞v����;���L���,��-
�"g'd-�˗"����/��.�q�]´�q��^@��3GF�LB���Ε��;UI(52��1����)���O���#
�lq�Q�c�3��D:|�?���ם�[���N�&����Z�c��|#5q���� ������e^k�����|�o��]����~��9�,��6��/��KuhG`م�Q9��6���fQsӛ�L�ht]C�q3Ӗ��Z�M�G��J���H��El�D
ɤ�)<u6�E\'�[�S�>;�8���?Y�$�<���PA�ֿ�c&<Q�M�cl9��XA*�`��5���kR�`�0;���V�giv��@�H���k��6����TI1M���/��@�Di� 1��qĨL�7�͏c>zirfF�U�cP	�ٜ�:��2���:=�Y�K�3� mJG�S�`����C �@8O��8M3-kD缒}���t\�P?�J��z�З&7��a��x���䪛[�Ebp�D��y�D�3��EȋS3l5�e��G�q4����w^ ^2=J F|e}�h:��wzɣ��F��tL��&<� ��Q�3a& I��$�]]�r7Fl̢�����)�(�(����0�N�K��B@5���_F�M�d.�|*9�x����S�^D�zA�*;L���S�Y��O?�������|L�C3䚝��{9��P�O���:$P�H!gL�zӸI���!���J�� �w�)X�n4{#fs.n�G��6���N�@(���U�iX�eӵ��Z)X�8��H�|e)������ݍ��14:���O�l?�y蜥�?����E��=L����`��K��m>X�S��i��G��.KǗ��U��<�f���9�2�Z��F��Lʖ���ЅN+w?����voP���Bˈ��N}�ǜ�M��
�QA���{,h����$1۫nA�!�!� 1��/ �����x02�*����d�l��c˦�a��)���DT���zm�!�y�o���5
��|����VM��M��*�C�}�{e�sz�}�p����!;�Jb\
��pDGFs]^��D�@��.�@��DG�Z��H�; G!HN��((������)���X~�k��{���Bd��4�Ȁ��X�J c��D��r�8��3���tћ
/�1��@K���V��x�o�!^���hh��$&�Y��S��NT��,*k�K�/F.�y=0�&��<��J���h�􈻐	���nR83�֨��"��X�?���0![ 	p�q�pg�/�2OZJ�6`&�Z0�[+h�k�9�;p�r-��C��w�wwc_ys��EW�NW��@e�q���i1�e������p�,�p��8���Z{���O��P�ֆ'P�m<r�ɗ��4��̾������}�Fϯ��7r
�N��>䶬 !�ѝh?�5��X	����20��o�	@�8"j�w�V6@yEc�F
^ R-U�G�/tq���Uϭ�D��p���9m��w�Q��m��Bƾ��Ǒ�I�q o��m�944L���ZPɹ�c���}s3�%`�g��Q��ȋ�;J�;�ފ�V�\�%��0��7A:T�)��M��TN�����Kc��!.a��-��x9���q:;Rɴ�UE��>�4�n�BD &(h��H7��W˗�$��9w!���g=���J��:=���
rz���ڪ7�u�׽�u���ޘ����ٵ��GE��{�Bh� ><"�n�M�@�@L(��tJ�?��_�G�ux �h��>�Y��j�Vp�ii��hR�l�փ���>�
�$%O��Kз�4������<�� �U���,��.�?:.%�����j�X��;B��z7�ݞ�2xN�r��t��Qt��J@j`�F����i@�V��ׅH�+'�osS��<\T.-����Q29;aV@����ΥI�t���H���^��aa՚H�NF�Z�,NS��E�+�y �y�?�N���"����eI.������Ԟsh~v����b�dQ�Ltñ�n�?Wœ���K���=��|p��f#�h

���2_|9^;:F�1����Jr�k�)�i}���>mO|l��i@K�ۑ�{oA|���7V�9���s���B>x#U���ᆹTȀt���`ޢ��H��d��f[M+�Jͣ�Z�m��c Z-�-n�@�7R{����L�8,�F)�w������\���
�2`Գ���ue����Jv�ܿ�܇�/���S}⋖}w~��sC���r;J�0���f)|�؍	Y: H���K�:�Ѱ���/���rd9 =��&�m���A��j������r���ٱv��;�AZ�]r*[�������������|wy�/��.�5�7�C�b�2���B�	��ޅq
Y3`�?�>�
���Җ=�������5P������c��M��*�i��d� ;	Uӡ�h`8���׹3FG�M$p��	ƨ ��h"�t>�T�_�U{���K*]ׁ��c��gERy�.����Y�ڣQ�C�<T�H�Y�⠢	Uظ�N�Ǎ���J��O�6�e��L��:��G�'ư��q,�<9GZT/����kQQ�dBn�d8����i���J��￶F�#�S�'��!����+��>���O�b]Z�Ů9Uc�����I�kA�`����#	h� ��{*n:�d�N�k��7c��ӊޱ>��fVЦQބd'Å(i����O��b9�>0x�G�w����:J���Kղ������}������b{1�G�-�b�AĀ�OG����{�F˜�0}����Դ�-�?z�9Y&R�M��	��;8,���'��q��@���c�Q݌�Ն�b�@��'e[]\��nV?Ϯ���Nj@�b���j�]�����5k�/<J�r���$��*������Qe�e�k�yU�J�mb�?y]4�}��VhPBG���E��0���@�G_qpe��#Ĭ~�3p+Ȝu��<��a�R<@�M�j��y�ww�YИ����EPH*�l�Ԡ�Ou<�O"*ŋ�Ⓦ �r�Jؼg��]����?��T�6��C�'hImvv�|�a.����S��]fRꁆ�Az�J�R�O�k}��զF����F<|1^uϨ��V��m�}��,n����2�?�/�gK�AG��m��*�?�`�5*�f�O�G!	���lܭ$#eTˋ�띌�oB����f0&�Ȳ����C#��V�>��c��T3��vU��^OSL��,7�S��-˵�Q�>��pď�xr��?���	��,.�e�\	�9lGbN��9��)�c��/ 7y����ut�[�1�M �k�,�n���C>ˇ�7�U:5�@�2�ڠo��9 ����E%����� �=�sZ=�DA��D�Z��-�
x�rvj=C��I��-d���F'Z�MRz���Yl)�#O�AƏ��/W��ul�X�:a�<B��IW�Q���o��~~�zr�gO,�+�O��:/���;a�zuc�_:*0��H7�m�E���D,D��)��?|�%R�Z�\��%t��{}{D�$����k�j���̉����nP��u�9�t�BU�$�t�d�z0�βҾ,�&>�mV���>��,3f�b0U23*3��<*����u:�u�&`!�ys+���:�^�1>6U��l(�k�FZ�+�����y�5.)��e�Jb�9�B6�t��~�z�j{nG�l��]�"�Ǉ/���f��Ê�A٬j �z���4�f���C��N���*n����~�ZG�Y/�~��088$����D��B;!WT�u�/��`��$
�0��o�����̉�9���=��n�>�q-�u�
0�D�$��o<���� ə!�?��;�5�*�h%��hU�s��[�*�������݃�'Pi�ږ��yU:��LO�m��g�`˅fG�z��cx�R-m5�a�nI��S"��#��S���"�-m9����_e�Մ�f������,Q���7�G�� ���}t��J:_%��x��z!�<��,gF��Ux6���t�� �`�r��q�(د��g�:�����|+&���%m������B�R2Q�t��;n�������D/�/Y�Tƨ������?ҧ�W�fN�l��J�G��[WX�`�:�V�f쉂��<�P��� %Y,����S���Ѯ�n���D͵bD� �BS���y�k�H`6�ۡ�(@;;�pW�k�jq����i�F�;�9�:� ����E@:Q��+�rOF�� k9E������.9J��!ZGLq��!;�NŪB·�v�Ѻ �Uʹ5��n/Y�?4W#ء��Q�T��\��}��S,��W|7�R&�IX퀲Y�O1v�	����U}��h���)Oςͧ�e�b��6���@)�C`���$W���i�����|���F��vP���N{Yq�{q�`<�q9�F��ѥ�Gh�$'�����ͦ1@~q}<Ly�6ŌqT�p	e�_�q��,�g���w�H-� 4Ҕ�W����[C,"��&�]���B����aj�%��w��|ٍ�{��Hyv���b��L�=�i��U�~l�"a8ؗ���Mƨ���ǁ���[8���j�yZ�%�������_	 .���I�cy���'&h�h3��ȼmi��JNt?�o�'��tq��OҎ�@�O���B��$���"n�|7�=�-�����G�v�9} ����-`�kaQ$�̹:��_*�.1V�}|�۾ϖ���0�6®���,|���]B�m�V���=vƩ>�;).r�(�,c�j0d�d�u�n�k��w/n���o�"�Ғ3��3H����/_4�e�J=��Xg����Q����^�s1��`��P�����3�u�lf��p�ʊ_+F[����C%��A�g�| \OC�B7"�ьН'��A���$o��ޯ�->MJP�O*��J*l�ʎ�q`4��y�pu��޳�����"�":��@�H��s�����X�?�l�.���w�g�++�(��`��A��,sl9Q�D���n�9��%!mto�b ��X��BV�q���Q�c�-6�NxͶ�T
����Uz�� ���W�J
2.���(��`uPs+�*�ho�V�x)�]}������F�ƁEI�y{�F�ܣt��V����w �6n�코��I8���tV!I$2�P�*�НayGS%����]q$,�}[���i�j� �m���[l�{[�b����(QfA�%u]�'Pp�A>d���0�Z󯡭��Z������}g�G��-���b�I��殧*{�G� �iJ��ͭ��"E�ʫ�!`w/mG��	����`60Y. VQM�D�����z��'xD�;N���!�>��F�qX8GIm�o9���uL����U�M�Ih�n�V���r�� �(*���nG����[��j��{�p�J:䠭)�:r�i�BD}
&΃@R��<�"Vn0�2�9;�c���ڊq��G��%v�-S̩e�ds�]ڈ����Rیm�jP�H�x���h `dX���:` ���/��ro+��'��GğJ24����_>���5ѡ[m����lҙ��1�ꙥ/%*�a�4@f��o-�n�Ū#�3A��D��YB��%pr���,e��h9���F���̥anHXH� �w{,.�� �����P_������e�ը�z
��m��d5�Z)�bht�w���G#�!��hR%!��ެ/^�0��iD��a}V��B��o�n����(�x�?d�՞����R���UӨW�׈�F�Av���D�]+�1�b!��Ji7�
���|��"E�g�R�6���wpd�ҵ"a9���़��Aгpp(��ϣ��a*L�{s��\���4xvU�~��S-�(�4Ԫu��Q����xh/)e��H'xmZ�@fW�xl�D�b��1��e50���`)B	�*_��$��ݽ�6�Ƭ:,hQa7b�
d�n*�݁��x�����8�~c��U�o�7�;牮$�!<�N���T��>��B�c��K�1
��9�+�L�]6����,�q��m��^�F��]�{6�MX��pz��۫q�g l����@=�k4��������ak��G�*���_];};���
���9��� ���UOA1�Bwt�G2��$.�)��W�]����o��X3�W(� �*}�A'��.��DP��;��s��~�/�����X��~�F(��V4�=�6���<�	��5�XKq`��֨�X�^~��.&M~�_�=�Ġ;���f��
`�.#^N��(؇�YL#&�6~�2�nJ��,-���ʽ�H��Ք	�b$�KX5G�C�����jzψ1�����Xq�)��>�7�qF�0��Q �'un߹#JT��B>�w�n���֙v��w�ͻ�z������� ��M}�|����K�Q򘫈Й�;6.I䵽'�'���S! Lu>�Ե�Qk�$#;��C���	�]Z��=��,��f����s��\��K7*��pjE�uU^*�h��5�fyW��WCЁ�k6�"�xX*>�J����\g�e+��x���+�.p��>�]fm>e�Q>26�l�27D /{��G�x���%2�����LН�O��b��G,8�R, 4�qN�pI�K���W��0�* 
� �75��_�9+��pr�7��5Ϛ����]ĊX.A\W��]G�^]jC]����d����0�P��"��F��κ��D!@����A�.J�6�۴� b�ȴ��g��ǽ�Rn���C�K��?�2y^���)s�L�9-��*�yj��@8{M�C`9a1.ť����o~�6�s��uu���\(���țߤ�*b�2��A�r�Z<�CA����Y��
N������(�8����ҡ�8OD���%������ż�	�a�d֏ْ���e�~K�7����WSF�M	眺�DK	�p��K���y+>�EӗP�H�|�In2�$�![XC�ⶻ�!���%���c�˥��� ʷ�t/j��f�w��tY9�����A�6��#�߃��q��s�qm�6TpLb�>ŝG��^T������&�f|�k�[ߪI�%�E���_d~�A>[e�e�h��E����GB�GeRg�����2��>?��t��2����ip>��)�FZ�Lj�at��n>1y�I���?K��Ӯh�%�ML{}�&+:i���LЬ���$�1\*�L���u;Y�_��v$z�ێ� YT�#��b/s��ٞ:d��FѐG"���L����M����η��,U-J��V艻1�N�����3�"�wĂ��^���U��ޓ���R�	�T���/�HD:Ƀ�����7���:��ϵ	���u�7B�����Q�� Ga��V8z�ȏ�k�
���_�@�v3m#/n��;�l�����Z�֔�rA��-�8110޴��R��
y��A�jx��e-��轑�Σ.$���&�H��PY���Z��d�n�>�]��A4��"W��%/�>���{i���_��6�&~8�'���nZ��+G�0/*�����H(��"�5.�(]#�i�b���8��k5��G(�S����V����M��D=�N�_#��.k�C���V����#�����fZ&`���}=Y����XP�C�5�����f����s�����;�Q�M�� 	2r
N,Y	���;�[l������
���<���w8�kE;���kW��w`��k����EW��4M�xH���%Q��˥��[#�%��\�n�/�YN������)��Ĝ@0���ekg!����|C>ŵ��g\�{�x��ǔX�.d���-�p������(����J~�<����c��/�X��M�KA��Q5�=".L��'j�y_��\yPDU1�9]�,虒�lq��j�D����l�M>�^v�
� o���9�~kfp�<��!�L��?� ������L�U\/���W-���vIpq������ȥ���f����Y���1k�� ���B'��L�Ŷ�l�
y�u�y��u��;��<���$2瘍�0.&��H� "UzXJ:�Yw���1Ӫ�X%��[]�I��k;�p&L�#��#�~��1�
���Vw�X��a[��w2�P A�]�K�����8Y����(E�����;�F�[ �mxG�៳R�H�C���5����K�X����(�Ԍ�zN$#/T�&qe�%&V薠��K�̓$��r˰,�lW���Jp� ܧ��u�*�9�nԷ�����j<	���O����ϑ������;�|�3������Y�:B���3��x�i7|���V<����p,����Q@~��J����g��:?ZWwK��?A��o<��m��b{�-c8�&2�ac�Ú���kޥ�#�g5��lg_�I���N���]�,-fԫ��͈`�˖5���x�lΥ$��%3Ƀ���}��|y�h�3�2�8��ţ���5P�6��*�K,b,�U�~��<۷UG�<E����G��S8^��j������d˒B��\�?�*�I0���s����k�����&s�.CN�7���ި��A�3pˋ��Q��S�óB�@ıV䵇M8����D��RM�t!X��h?mf:h����}=�7~ލ��W���@��R]��t^�lzZ����y���`|�k�w��P2v���-��ګ�+��t�%�X@���c[�)*L*�Z��`w4�k<M�/	�P\T��}_:ᑬ�I1x�����.{�3I�{�-�TT���cfw�w�5�z5�����/ƔUm�o��@���s�R���ĭ}�pk��9:�V���<�V#^��lҲq��Cy���������݂75^����GDuYӥ6���ً2�ʠs��e/�ˠ%{T~�ɳa��=h[Z�T���Cq$����96��Q��U�af?���+����V�Z�\m95�����G�[j�R�'�����xҴb]��?I0˭_O؉���f��]�M�:h��~���م�bӷ��EB3!�}+�E$��"�F@3^[9����Ə�Yֿ�<��j@�0@28$Å�,I������Qb�֬,��%K83�m<�17��z��.Hբ�7��oePՆ8���i�ҖFv�d�}߳RNlh�f�%4DG�_�lћ"a)�p�$TLK���=�(��cƇ�N#�̊��!snN������R��d�qB���Wr�ʇIi%��T1��F.�e�#*��y�����������?ҿ���?���J�s��� 娂����B���9��Z|���q�0�_�?��u�h�q�޲������E��Q��埃���-�w耫��5�[9ig��`��ʫ����b�8
&��	��*���;�"��V��?ư�n�QK�2�-�#|Z�Ɲ�G!u{��Y��C��)pDeE����a/����<�O(�h3!_�k�;ydq�����Z�w����w%3���ռ��ضB%vO���	�J�F
1Om�\���L#4"�x��Z1�9��@�F�3L�d�W�ղn�}މ=�&��O�џǚ�l�m/au!�1��}57bǎ�� �Fb��R�3I�����J�C�N��=_��ϑ��i������"H&ߋm7�E%켾�SL��� �����J�@����|�	S��;�K4�
��ރc��+�2�ZW!M�M���)���2\/s�vH�e��+��_NF��t�|����L�gҧ�	&Ϝ�jX���R:�sNPk��+�A�<<ש�?��:�T,|�#lp��'��ZFwq%�$?{(n��^�����kDOG����E�����O�A	o�
2�o���5�+�"��$4�Ѵr�AW^А�d��������~�\�*��Qf�vE����kc��=�����+<!N��Q4Ҿ����	m0�i�LA��B:�]�P�<������[}eRs��b�]���������/ȋWƅ/��kX��:W��ŉ�
c����Osu������J����H�zot�]k�c���ň��;t�V���sK!6�3��,����F�V�D��IU�����˃��̡�5B����3����'m�Ps�DXr��;;��}��aI�fn�ar�FE�����JiA�w_�:@�����J�FxGr�.(�����%t
01�������I����G��E�g��X<α_>��˺�����`H��p�if���F
t/����V�I������є�;��=�~a�[�% 
J ��^pE�H݈m�2s�uo�O�g7*ڳz��6�}�#Q������l��]�_1��w�]�&�υp��>�N���%�ϥ�{tJ$��k�uu(�p��xH�FŠ�C�C��`yU���;���V���L�+)�j�����fS��I����\�4����b�[�h�0Pu�R`|S�Hy��xw��W��H�r�UO=]��9�����8�׉Q{;��#/�"��)��K�(�>5d��]�lHhC�?��t�7~n�������6�[��yp[_�?��C�M{]�
߭#�
hn�,�Υ���!ؼ���;j��x�:ؐy��gݝ�i���a�_��,ci��#r �GZ�U�<��CI�3��l�����S���U��{��~�2r�nE�Eiu��U�~-e���#Ճ�z��Ǘ*�I��.��<9����y�Ώ��}�j���] �qCy�����:�N20R
IY��6�0l���)����;�����v&�4Sq�;'�#��A!�g�T�`�g�qp�R��o�/5�W6�x ���|	ICz�:�O���W�8Z��.U4JO�^@��l��[$���hO�ڋ�y���z:<��f}���L������C݃�Kۻ�M�?�	(Кz_�[��X��I�4+�RϺX��r�@�cB�eɒ٢�$�k/H���C�FSK��)-������J�;Zf�mk<:�� U,n�>H�~,l��7ks���&Dk�H�/ `τ�|�܂�<%�]�����^i�n&�i�8<�Ź��'0�����e&O���ʇN%�|��8����sF�q��/�o�F�L���6C�e�x���hnBdd0��i�_����U�6F���?�ڢ�1�Zے�g�2����d2�
��.g���D����A�on� �{*�H��,��?�ݿ�bf�"�cE����{x�����X���2`�7��X���+�~?�A��(ݱRI����cz�B�~���ϼ3׌ZQ;K����~�A�gM#1{�b�ƥA��U�eWٻ�ق��QƁ�2Oο���%��V��u-Ӧ+� ����nzN�C���7����b����,*�mX���-��Wy���渽�Ic�.IF1�Ԕ�6ڕ=�����h9б3�(ĺW�d���H��� �W#+��D��.�ӦŇ������І��h����L�63/�B�A�c(A�Xs��F�(�?����Ś7d˅c4��4�4-n�H&9������D$�
BƎ����\�g�9���覻����?d��rdJ��E�{f?b��Я��z,�w��R�<�B\@x)��_�I)F��͠��ʄ)����~w�P�;�=갧aUVX�Aџ}'��]F����t�����"^��n6���A��a�87 �J[��
,�5N�OG�u����wN��O؛�n���Ѿ�� v��c��g>��Y�/���׭-<��4|�;!���N2��u}���C!x��s����^�j����� �P���f{Sެ���I�V��{A�Te���{"�ܷGr�_��%J,��:���W���r�v
>�dZ�"�;��;�򂮎�އ���9,����I�96��6��w�I��׋�R����#�s�e ~%mS�6%P,Q�G��3�%k|^h�h'N5ő�G�W�@O� ���ᤶ(g?}��d鄯�uY��`3�X��?�"W��ubfh�Y�ٞ�E������x�1�*`]R�9'L�(������?dI�eC�,$�.Z9�C���.�&*g}F`�?@��l1���Zt߱�M�!�)*qY���,����si�!�A��ݪ��TP�d�q!�b�ۿtVB�aheKV�
 G�m�P'���c�yR�i���e�u�ʞֵj3�n�-��aC1Q��9�8�T��).�Κ�c���|m,Zp�-��Q����t<z��#��mU{x ��8ķYjvc�`R�W�Í-~�~�U�k������KmO}M�
la^���V|�r����ԩ����B.�"?���t��f��ä�ǘC����UlBʪ��װ��)�>��`��ˍ9�}?6 9W'����r�M���V�'������Bk��'�<�G��x�b�2A�������0݈=�A��]��D���/^�O�����;�7�$n�>}��`�I��01,�(($6�����'�{6q�V_�ܹOz�*�e��P�?��AL{|@��va�!DB*��~5�-n;+j#���^���]�����5pcHc�,T�OR=�}0|'���ˀ�CNxK`�Ϭc���P�ޅL=pR�7/ w���c�5A �F]����Q�L��m�\ل����Z���2��J睬욺c���rX�sEKe$��\hR��~����4��5��g����Iy�LB�	fL�-�3�T㏵z�*��]0�q_v*,썺p��<14�&WW�TN����lxcq�~��m�E�����o䉁��sR�E�L�In����`ڽ{��/�>M��ĶBCւ#�����GK��mI�X���C瞺�|�������&_�\��mA#P��&�k�d�<q,ws����!<Zs�*ꂑ�����p�&�Ӡl���d�i��H���H��-�%H�b{ ��R8���UU��	a_��k~F!��u������a���#�@ݑ8$f�:�lRaZm���X]�/�����1�{!W��p�v��o0���'p,�D�X���[PS��0���*��E2�Z��� �2�F��=�V������3��Hfut��q��2P��H���z��=Uv��1��!љ!�iNf�:A����mCfoDb�Q�Ol�+D��.b�ߜ��_����BPtq�BK�����=�"(�g�w8�����8cn3�`�����ST�,����B9V�h�V�}~w�`X�j� ���L)�_qr���\$�q'	�H/���bE4�V�'?��<@9M���	.���.��5�ĆH��WQ��w91aSI�tk?Ƅ&���#D���?|��	m;J��+Qw�b����+��&R7��H��	���6(\�tK���
���$S����^�}���(��ۯ�Jb��˸��m9���^bԩ���񋟵c���A��Q�Z32�.��
�pЙ��F� �`��d/��z�]R��Y�'����}^�g�x�4��*ә�.�Y�CF9"a�X���Ӑ�ȺoIz߾S��f/����?�՜�����O�I��D�V���b��B�n]����>#�|�����㜅���.�d������~θ�%|�Ȗ��7�`��J,�����Ǩ��Ӗ�}s���0�힄���dP<��2�'qZ�,����Ni|>�g)H����%"��ğ�%����«������H����S`1���-��]�j���t�%�F���S��<PB�����=��u_�8�s"s�l4q�����ۘz�_�m���Д4�9�&�A1<ɗ�(G�.�j�S��Ͷ<�}��%���o1�#�]>�kM��mt��F;��ɇ~?#vW��CuE�\i�:���e�Z��xS����&�Z����Y�d�
�7ɹS�w~���-CU�ߡa������5���ޏk[
�al�Y�y-�Zw��xc4|�=�OVk5]1:��C�sJ̅�D�\���[^��������UV��&�:��"�&(����v�2e"��Kyo��]r�Q�G�$	v625�M �zV��#�3�%~-��R�/�].(�t��+x���bW��?.�=?�J�4+���wƺ/�:���nv�c9���)9���1���+[G���)
���*�ﯦ`�$YC���
C�b���@<qT�2��x���5����8�k�BR�в�s5�a�xR�44��z��X�x��w��?�9/Mmi�#2o���:?(вp��䶷Ő�9��J��E�*���2��Q@�u����s��$t�i�'@�(q��5/҃��b�es�fK��^���K�1�Ē�I�o4B��W�@����b���_�ӷ�6o4z#�,�����o� <\�0G�O&Py��C��TpU�H�}p�R�����	��L[�X�W�2��'ߏ���s��@c� �����K��W�R���*��h%��ؒ����+�V+n����,�+�3�	���GmǬ������.�̓l��&��}q�M�?G ����h���,9w��g�L�C�k��݁�jb[y{*8���nKD�1�#6"5����X>�y�6$�K�I ֓�LR��{��ð*��dN�M�,��㇡�qx3<���FT��%��*�Y_Lб���"�v�(�.���if֡308�
�����v�o�<_9�ՙ&�|a�Bwq����/$)���l�.�g!�h:x�Y?��sW��ǖ�¨r� �g�7� ���zߝ�i��,i{�ֳ.DY���)sJ�@��@�u�d�q�wV��m�����J*0U.V.��>sa7ɤ��ə̄35zJj���Q�6���Y�k��~�2�j9��5��F���%H�.���_ ���3>���C��;-Z��ѬL�,�͠���ƌ��v~`�W��ҟ�pH����#��f਍�\cD�װB[��JD���[[�1:@b#����br�=}�
V���oǴel�x�$"�w~���+�����_���eΜ��-�0e�����XZ:�����^��^ZAyùy��&�/q9�*(�%����c���4�g[�bj�3$����.z'���d���O�4H�p�iv�]ϣ����oҔ�?�#��gg�w����Z�ј���`J�Tʷ@S��嶪���L��Ac�h�/Id�ҎP�YT���J�9�Su@�����8G~'�>��w��%z��@��������/��W���Dw�!�<���}q�A����_���+���e�K�<s~,Po�j�4UU���D���i�A���c�&T)qx��2,m+�	?�)�,{u�5�4�<d"��R����x��6�d\�z.��g��\��u�<����e�X�)I�d^�O@A�߂ܰ/U,����O�yCF{���<(���ԈvH
���F`�s[�w�O��,,�M=� ��:�I���0^��R`��9�U{~�א�mi�*jm����5��f�F����S��O]�G���<�[k��_�K�a��zݺO?�1~�d�cm���Z(��F6�⾨u��"*lU.�O����ѹw?��������4�:���'���;�������t�^}��ng�9���抺"&z���M�^�!EK)����s5-�\{�)H��{(�bϥ���������;��>[M��ׅ]��]��&��ݠ �J�
W����b��B�q�Zb���m<�tkS�^�E�eנ��!�H7�����x�C#*�󱇨*7�[����?i�L�
.
+���j���Up�&�ar~ZI��m^��	�a9/ SӆpXuE�w7��&�H�|D�
2x=(t�o��T����	\�,��x6��2lz1�jZ��]���X~Z�)�!�:af)�ɵ؃�Ϋ���Ju�.��f~j�O	|!���kx�����b�eG�W��A����mAo�I�b����2=���o�������Y���O��c˫`�<t��x��Hť�2g��z�5XI�V�����O�{�/ȟ��¸��U*�#A�*Z���-�v����e���m��+W�m�dQ�i돷�=�3�}�((?��ao��DUePƞ����G?/�e#��"<�xP[��u��[$��&��ݺ�䎨B��Q|�,�X��z�]g�z�4*M��ѷ����6��+;���~�U�oX�(�ۙ�!Y׺�~fx�K��/�85�����Ӥ3������;���0ז��O�"^�$K��=]M�+�u��\4�;�����'q���/,M�<g�/j�����>����6LK�X!�?�:�}N�jҜ��&i˗�i��X�kCWs��giʬ�NN��ڙӣ�O�V�_|U ��:t�j�SI$��9ア�y�i�eBX�!(��4H�RpT�b���b� [Ԩ5b5��r8:���\�s�]q:x��˴(k���F����׬���P�4���;i_�VKCJ�q�t/�	Zbz����K^����&�#�� 4�Nyr�h�B#z�f�Z�~E�n{��5�K3��`�r�	E�E�L�]1�;Z����"�CtI���P�L�sP���&1�}�;�5e���"�L=lĈh��������`�IiBM旓�%mqX@>�����S���!�g"��'��C�1��m��¨Oŀ�%��c ��3�P�ͳ�څ�\;��^���+РK Nݹ�'8\���@8ދ��.�2��M��d�É��?�Ԅp���m�C$w�1\P��{���(:r�`����o:IA�c�:s�gM6.Cz�e�v����m蜎��%���nF?-} 3#W�&YFl�����'
�#��%��5zOq/c�ӷ%o[����>ẓ	�Y��.(�6�hn+El�R��U�e�h�
�i-����L-�WWs�}���U�0����)i�L�p�xS1�7.Ű���[=��Jvo����T�� w������L{���gg^���cyS:��:����4h�������q�$x��5��}48�hHA�7(�Lo�
���Z(輨U��d�G;��xs\R̚�E���_T@/O�I�������:=��J[�؈ �|�0��
��W���./���ǻ�V�ى�LC&�T��5^��0W���^�����Nȧ3�0�<�n`�0,{y����"�)X�L�0S-Ɲ�2]��,���d�7 pESJ�d�������egH�'o;�F�A�:���@1��SjԼ��u���@XMȂ+��TM.m�������,���+��n*f�\V �'�X<�_O���ݠ�eg����q������&���n԰0Ҋ%��I�^l��E/>�h��#gu�!U+��yjo�F��F�����L|��<p0Eo&�;�oβW��~�=*��{P��M�l ����L���%����
5�H���t ����p��oN�~!@����g�&5����ym��^��P}�AJУYCX��ZF�X�+��Bc��ܙ��5�ꎧ%~a:d׈=�4s̍P`��]��Y;��h���n��Vb-����%a��l�~<���ť��_��L�diBa{���寘����<�,��:�M�{.�����!V˅#��jƚ��W'��BA���8���ͥ�Æy��Ǭ�֋nQ������Ld���p�}Vv���u淮�`2�gy�c��S�@1���`�)����\��X'�:-����ڑh��$�]����V�:ܒnq��k��VS���)a��q��ۮ��H���Y𚫅�X��̇]ˢ|��鼀�+�����z�K"�������L�����8����D7D
߷��쯝xg�8��_BC�k���p��y�n�����<��&@qe��O��0�zb���#P�ٗ���R����?�%�gM<�L2#��eY i�+	]0�%7+��f r�����NJQ����%�\om�S�Fp��b� �20�D���P��u&����_Zh��o�C��)��>�~wM`��g6Jb���h�M��a�lK��ذ���
�r.���x���d�������r����^�VЗb����M��G�p���&��oq6���$�)����j� w�:�@gMi�rPg^�L��lr_�8�װJ(�G�����{����a�Yj�oc'?̲�F�J\4�L���p}�XAp|zK�9.�/ )s����vI�(^'�4��OAM�vc�ZC4����ȃ�6���?48ڍ�Է�	N�&�{��e��p�&ub]�y�e�Nd��M����t���dd���64M�����͙HNz�84z*ne��$i��c����|��iRs9
vo�@��:x�Mot�ݸ\v3{5M���8AG��đ"<�w$��4�>J_!�!��lO)�~H�?}]sq�jᩔ�0�W�4k��v'�A�j^ʢ�f�(���~p��NfAwظ\�n�Y�{�DѬ�NXhk7�o�}����V��`�k��7���fb*���>'�'%�S֊M��Dg"�ꝕ!���.{4�����5�zx��z��}�oj�:$���@���6�?�軯ԭT;����d��<߇����t-���N�t/��*
��kY?!a=F��k"mH��&0"��r_>�ф�~r�pn>�j�B�zU�1��2-���*U���4�-����WU��X�둨�/��m`��5�[�Ƹ��fd�t݌��hAXؕ����̭U����ۗx����[�30�${��A�ڜ#ǈ|�4��陮�R�ڔo:.��k|�%���ۯ�CD'C,�[��GQ� �c���/�
mp��a�����=���q�ϳd3��ryH��a����Ŋ�.��|�D����2�m�׶.
���&I���*�#���2��gJ���A��7"�&�?2�TH��{�x�I���?j�w��ZO���|	G��)�?k*��yaҿP��9AӼ{�c�.eT��l8��[�j\�܏[�F\�%
����2B1)�E��8��ual����L�	�3�����	�/�i�&1���)�e�CF�*|2�O�{3���V�[���T�E>��B���[�sS�����M���7�q�*il�
�'�E�_PX��l�~��\�x��(������r�ݥX�I7 �"�,%��8KΜz����˞�/�@���#T^_!Ol;�k�Ol�զ��iHo_}��8�XQ�c�����D�)cNy�� ��c���G�ÿH}�����ɭ�d_�[�����`|�$��LϑyQ� ��	'JQ��\@�������4p�(���S�S�f�����l�׉쓝zb�払o�g6�����aH2T�T�c�f^497G�6ޛ �,����%e$ �(�6I��^+��~�"íw����@�ϓ��n~�����K'�����8f�ٽ�Mʲ��D!��^9���M�$�4rķ
s��yc�<b�n��Y�Cj��J]8�\�ό�Ny)=�_Ɣg!c�/v��J�yU�qִ�`d���X7�z�v�l~����M�T �	���Շۿm	nk��sy��;C`#H񜢨b�S\�A�C�Fޓv�����s��l�iO���L�v��Z��h8F}����]��D��̃%��U�+֦�P�
�t��\S����(���'b���TX,9�(&宏�ZHj�ܕ b:!Dp�\F���C�m�����To�H��m�ƛ�r�����7�$é�3�r�����iR#v4�϶?�I̍G�d��E�4L�4��*�0���J�}������ʘ}*3A[X8�=u�,/�&���@0��O��a�"HUC&���{��R�;�Z5�!��k3���<�6��鎑W�\��Z�D>W�黝��鮔� �2���fu��G��zy�}�.����