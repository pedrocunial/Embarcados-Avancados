��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�cЌE���MBvqN�-�	p�ЪHQ(@XiI���a��B�GH�_J��@�a�LM�
k+6�}S�x����)=t`�~3�z�p��_�������!��agZ�b��5���� 6
��b;Q7��*aPu��g�<>'4+��E0��Jޖ/$���Ѻ`��)�fH��0��k�E�.fN<!	e��Bۄ���S�l��Vr�-����t�o�=��B�+�-\1�W��OMj�N1�+��Q�hWb�6�ޱ�0�%И*� o��&�AN�e: �S`S�>��Q��_�3><QB����fA�������'3��uQ~��5!XJ�o�p�q��/�q��ɻ.w�6g(�u�ɲ�Rmfφ�i��vz������m*��[~Xg���&����X�p7��>�;U@8������o�~��������^��.�����҅�o=@�Fb�jW ���Jҳ�=�^m-���K��11i��f���S�Z�2����#2�'�w����u�FeA�ƃ�B�NC�&�}oW���O��LOa$��｣�ᤝ�|��p����51+z�R��4��#OR��b�n\��Z	 L��C�҆�6�"�ΰ�v_]��X1�U5�V�c!�h3�x�O��h��{���<�%,�j!+D�4��	�4ID��~��C�\�ؾ�� `?b��lB��Bǆ�{�x(�t�����H
Snʇ�(����8X3�������E��B{Ќ^��(��E���%�޾�P�����d
�<�>B؋�g�:z7}��1�ّL�+}�7�wV��?1��V'VZUx��]�gO[�:ŽR� ��#�y�0z��^83�ᬗv\��j�%��������d]Ȧ��t4)˼� �H ùN5��{�Me�$�!��jY��M_��[L�k	���h� C&��g��� L��é4�Q��삟�б����Q����L�Q�\?�x$��ķ�D9Yy�6,5Xd�>���������{iU�~��bg��W�;#�c1���+�n$�O/�RJQe7G�,lcڊ�?�N�u<bX�Q)����V��0~j-x�+������v�pVVi�����`��#�>VY�ɶ���G�h���:9���������/a?&���V�5/�+�& ?��U�pA&/�G��Y\?��z�]y'�/E�ԈN�a�j�����JY����Y2�Q�'���pV�d7q1,[zO�_r�rU��T'V�&	�"��W�U���e�Zְ:<tfp1a��z�X[�N�O��D�g�s���C�-\'��!����^�ɛf��6k�|<�W����le����6�E�|���T+�1��?�.Hm'0����<� �'u�@��R��h��	�CA�MGE��Ap5�1�Jk��a�xc�5ʻ�7^-�Ґ���H��V��K�����lt�X���OP��Z��jf�J��3k���5�l*�fj�51b�j�|�,���U?d�d��m��ٵ�SM�1¨u/F����rU��v��@˭�o��Ȗ��͙���e�d�E}X����-+�n�s���/�|r�$-� �����j�V�O��#���bK�)J��i2�`����Qg�Z:�W�#YY�v���%���e3F�I���f�Zk_ˢ��j�CzI���H�݁96>Z��ϭ.�6	�}�6Tڱ���wG��C��Dw<(~�r� 6��P|��僞x|N��!8�����mt���K���=��=j.�'��B0�0xM��HhA���w>�ۊ�П�b�Ii�8P��g��Ʋ�v{�'�/��t�P2��uvYY�T����%�*�O�&cARO�1v���S�PZz����#Y�P�)�aV�퓱�l9���i@C��e��k<���H�+��*�R� ���D���"�6��Ņ!�b��;�2#>eO#&J��\�ז�A��O��/�C��3����Rp]���T�	)4�a�r
I���@���M�z0ԻG��5A�)���7��Q�O�u�"x���%�?�,r\��J,�?������<�hF�o����N�Oe��jŷ�+�:��n�/��1�@w+.T��Bg��:�G��0�D1�.�S {�۰q\biM�DvK�9��s%W��̑��/DY5`!�@��<op�	niAï����?7���#��u`̯DE1�C�CA��{��!n�S�ŝeJ�+��F芨kv&��^�;�'k��N�_ur�\�Q2a�L\!��G��D����3�����y�aj����� ��K�Ӛ��P[a���;hdĸ�9�<~��� �0�5۪����H�?�*��[������k*�RFO�;:IǾ��