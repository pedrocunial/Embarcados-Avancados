��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c���ѢǓ2�Su���;G�͘o� ����$�ALd��9��,ݝۧ�R���X��wP��1���p:�ǆ���]���Ļn��=�F�����W����O�7~�ֿI�ST�P��~�(��S����pn#��Y��PQb�,;�X�1Fq���Ռ@3���%�[1XU2)`�ս�@@��ܦvzZ˱��O�:O̽���s��۰1����0m尒�v�:r��4�,Q��J�ER�`f5y)�M�^��X�Vo�E��kO�
h�K�o�f��M1n���!uBi�%D_c�l�
��V�ed��m�V�ǁ4T�c?L�EtC�g-�����h�GnCm��%��@��s���_/{?�!{'�.����i�򬨓�m���ꓢ+�=�5
нM�":(�s;"�R��x�*�{�2%4 8!T�mzp^K���8s�,|
�
43��<-o�>�*xC�^yu_c�������z/�	����`.}d�D��_2Ё"a.x�	��'���� ��y9W�A�8�]홦rԽ����*/��w���N���M2	1s1>��(�����s}�V�-���@�>{<Qݶ6&�F��^ɨ"�/[x}d&u���6��-�FC�Ԇ,geba�E����Ѝ�'œ��$��7��|��s���ϖ�~�UL(��#9�4���=����d���6ռ�$�PG|��ű�Q���:�������b3MB4ĵZ��.�����=��%���G���Q��9LEN?%G���Y�f:
r�xC.7F�m�g�_0�t�Mf
�Q�a��L�~�4x ���#��궹�1f��'G
�	՛�T����} F2C+�ᎆ�����X�2��c��Yp���l����~�j]��m��`?�;tY�tQm���n۝lWT$c�`���s}t���{�q8��Z����?�2]*�������.[Z�����`����(���T=��O���"̆&��V��QS�o"}mB����h� z^>|L�?�;Xq:}�7)�g8�}�imE��Z����4w���{`�2ު]�t��2�Sށ�R���ȶt�P�&EJ7l�UR�e�9z��q���P�$�m�0��3|�X��%������&��̜o���A���r+�j�e��uf��)0,2F"�Y��	�:�_�6��,�q�Z��X�݃߀m	������">�-�#s3�NT�w��W�TIk<� �y�&5�Jgyo
��j���uS�\�v0���g���v�^%������ҳE�D)�v�j���ټ4�S�i?�c���y������a���/^�Ws	��+��>�9� ��j	Ʈ|�����<G���7eO����^���8e|�l�4����L6y����ɐ@x�ۍzO�{e�PA�k��_�L�8PѾ��n���������.1�kjָiL��r����'�)T�u����)ӽ�j������
��d�fkX<�J�)����:��uҔ� e��%-�;�J-Pi���^#s[d�{��c.�|P^Op�E��[
�k����--�bA,rkh�dw�k�ݻ��M����f-�M/�M��<o��{q��a+��.re���so���|�E�5�.����NG$Jce���;��4�y��҇D�Hj��p@�2c��J�� ְ�y\y���~~���?�2����P �MV�h�Z����~n��(�;q��4���2Ӯ���\�AX��@��x�_�/��e�S�Tp�[J����i[@�f��T2!Z=��~[a��L�6S�Xi����F�̜G�iW�)1�¬��Vj�MwY 76k�Twu�<��'>�@�܅锹��������D���VTC:k������sb��6��#Ƒ�N5�#uȬ�X]�	�<�r0��hf��o�ơ(1,�[w�����X�Ӯ���!��G��T�KImv��l�ةv�����ra�ϝ������z3���܉rϴg��-mb��2&PA3:J��r}���\����)�DB��cmV]�%�\*I���d`�� �U��C�K�QF`}����*.Gd�����"��=j$_�$��/k
�G�V�C��'��M���\�0�_�]���aA��L	%\�l��-(���1�yk��h'@��b�1�3_���'���WF0(�G�5*I��{�ܜKNx��߽8?����,vmԎ��Ġ˲*���Jd9E�����p��>�
:|G4�y7x_,��0���[���?:���E�|��)F���]��4��~�������8�+4_�V�4�����h��x-/`e30�P+���E���R��[B7}9�'!���A$��V-Z�ǩ�Tj|;��#�<�.jE�Wx��Eҍ�'���k��~!p`�	�0���s�g���m�W�.*�%��zUbڪl�����������q�
��5:�����睩lV �ȡU9^JK��X%�  �$P	���)^A�C��7����u�:D?�4D�� �����!&Ъ����u�+W�!S�RN��cq���85u���	[WNľ2�j�����"��� ��jr�n��rɺ= 	��[�;r�xY@L���YHJ���l�h�IOX3Y�%�S��B�0��F���Q�u��:��u�f}b�d7�p�o\M�T�U���u8LڒbpN�K��~M5�����pv��j����m\�D��p���qFz��9���N#l��N�K�>N�e�\|��9k]R��g�c�'���.^4y����E�c����?
���xB���Ͷ�l�:>|k���e&�|X9�<�Z��hh"�~��W�O�I�"�����pu�*Ofs?D�&������|��L�e��4)=��cS����'Ҕ��g�l�]�Ŀ������6��Lx蠧�x�$N͇{��q�%���� �=�{�8�j�N����	ܢ�/9��PR'��(8dL��m��”�H���[_'!�R½b7��m��7����,G#B�-o6E`�?��J����JS����]"�L�F?�S��Q����ͣ*rs�����Ʋdd�2������@=��ca�����rV�l�)f6��FVR��a��n��x,hS:��J`��(ʹ���_~sYx{p���Y��!��Q���@�x��E*�{�%9�>5]kK�CK��i�񄙔ٳ��{����`����H�i��~=�{��.\�A� �\�ә�a�d���G�eC����n�3�hiVVIj�H�}�*ſm%���
0�*R�	�8���?�zF���$࠵y�׿ӵ�\�$e�w�RpQ��^������&`�.�Gu���(��v�sqR	�\ȗCe�Q�[���PHʯ{���1 ���%��xm�QI*�*�����t_-�!_��п���Us�R/����f]�޴`k-�K�m^>�<=�BT&���4��V=�lB��9����P)���F��7U#'��x؆ea�RH��y���jI���˗�>)r-��ԛ�5���rp�Ӳ۔�
����9��KbܲP4	|ئ�H
ByA�E.�~�5���e;Zw�I�O� �����0F�4d�~I$T*�H*�"��W!ߤ��\^�,1�tC���$���*+`1ypx����[���XF������/��V"
\������A]u,�0c��(�CI�6�-�� �� :�m�;h����"���(�V�\f��(W��w�f��C�;��gd�:�eu��\�ɝ4���^K���� �$�\�Y��BQC��V�q`{wtE��r�F!���j�$r��S�wA����RALP����a��K��tF ��`��!)ҕb$��9��~ ���j��g�,�H!��H�L��7=ǡh�mb{1G¿y��"lU�I�d�m�������U�;�+40�#�9�4alXɂF��X���UWJ�� A1�F1���r9���Z_�|��j!P��ԙ�ْ��{����eQ��Fk�*_�����HV�6le�.@��
�dE�W(2&#d�YL=��!ظwE�����f��zΘ�W�Ԓ�����n�(�-N^���Ԗ��Y�$��1Ů�,��^�gWPI/HO�V�H���r�T��.h�,_�ؾ	�v�w��A]�y#�����*�'�b"|,�g`� *�+ޜFj�$Ȝw���0� �Ư�kA��́0QFi�4B5��R߈���q+���u-���ٵ�H��G̎�Cmz�B�����[��o�;��/��^̚v2��L,R_�cv;ʮO`���A�n����|+�|���P�-��B��?���ҙ��9�Q��f�QR1��RúF�=v�4n=�ZRj�$W�Ľ�l�������}�1�ؼ䀃�4�'�D�m��%��f���1t����"fN����x��G�������gN�Ü�ϥ|��z�Ȓ�KҶ]S6�OeUJ���=��R��R�:2�Ϋ�d,k�k'�<��$�=S��:��:�t���^��F�H��Ǹ֕�5��G�Rl2Ъ��V�-j@pja�.C�	���{L.�sq�0g3�hۈ�P�⬷6$Њ�����L���K~
�RD�cΏGXƻ�rp����k�R�K ���-���KA��=t��Ii��y��h��B-��?|j��r��8x�H�)�JQy��`������Ȑ�݇*����Q���W�8����b͏�yMu�Sf������1�k��)J7J�;V���hN�d�c�^��k����a��yn�n����Υ
4, ��ga\=�{x���Fb�t�����+n>�~W�2ĭ��:�.�O�ŋl���s�/�ts�ER�R��°l�:�M��齨�`��z%b�^�f)�� Ԗ�U��lh+)I6ԿS�=�G�J��(�7�'#D�Z�>f�]�nk�k�6P@z^��`���o�ۄy�a�Ϫ���+9j�^��O��^:�2�aF�OhV�C?���U�����Lc$��2�������z���+��r��f�F������B���A�R�\Fv����6ur�?r��@�B��7�F�= t�Ms��%����R��S�j���_CN�7_6� �39>�XW�ʑ�x�s��`0$�Xj[�4�)�q-��*_;��9FZG��M�����S���eӸ��$^u_�V� kQ��ށ�I:��͑C�ѯ�w��k�R�	�y#��Y�(��`$5x	��y5���9-�Z ��#C�r����FeVCcS5�(��g��k�s���I�S��a yu��/�OGl	\
���\���0b$�ǉiB*gl�@�klO��5P�8�%�����b	ʓ���~�=]����v� 7�6���"���{�8P��h����Z	�s��_~��^��]>M�S�}�KA��7�����ޮD���)�C����4�+v�	�#�Q7��3�=]�����P?�'��x!�,�[(�8m\�#�(�32�@w	���S�59�n�I�H��완�'×v�B�"�V
ǯ��2V�n��������o�$vc	X}7{��E��[���	Xfe����%��3���XZ| ���\�G%,��R�k�`Ɛ��PD�I/x-�ə ��A�<���$��mT��u�c_��_�r�os�:�ݐ���L���.n��2Ɋ��N
�ݖr|̳����)e�f@!�h�A�˞f �e)F�i+c5[~&�ɇ��A⢵��+�v]0�)WFm��&e��D������ ��=�Ү-Tr@�*'����N�x-Qt��3vꋏ���ŷQ`��|"�ۇ{=)���0��pk�ռ�ݡ}����wPL���dGA�s���Jcܫ�K4�'���X��!�0^�vlM	�Ϩ�~j�,;n���	�n�Eؙ]��H���o� Z7����+y�+������a��_�C�=4�qH�K�ug�h$�QSi�꽂C�i�(�����׸V����5�q�n�N+\r:���"r�a��NSo{${W�8��Ͱ	������8��%�Qo{����4=��5w#\��m�[f	ϐ�ୣ�����x*�*���=�����7�;�l�����2��$��P+?��b��q������_��Ȍ&׈l�
zb�	BWUe����;�6J9��!��󈥩܏"EB4q�vv��8��l�G(�?��t`X>oĚ)�$@�_��b���&�LS뜿"��I�Y�i�!�����R�0\�L��g7!	� ����/�)@z��a�e�q�u$u��JiӅy\6�V����U#!�N�G�.�x˕�LA��ѫ�}dndn-Fp��'�Sځ�N�����>{Q�%V�w#�^~����٣���u�;(��z��v��q����I��y P=� ����&%��1�XTW�p>�qI�ggU���;�\]���,A"�miȋ:�c����F�a��3�q�ms~TG���i����%y���+lU�'�Ӕ��jUհ�w� ��QU�?Y�;ϙ�>�tq
����_��P���V��^	���*���?� oH�N�N9�;������e	�y�e���2K|�-'1ʤ�nւ�v��̫`����R�r���NO![�f��),���fJ2�9��5�CU�R��g�_p��DHV@M�&���Tvp؂T)�NE2�3e��X�_B1�#�}������v��SR�A�U�E�[��@���ϭ��+)$y�,�=���$��/�1a��^��-WѸ���%���!����o��.�T�����V�l(a�;����@I�aB�����Ev�Xc�RS%*�����A��^6�k�Em��?��1�6�z��p;qY�PMP����,v��(� ��q�X�D�~̲���c�7fNV�;�-'\�I�s�9f������S_��7�*� ��??���{w������CĄ�
��FR��ơ) !��^}e�`%Z��]���dj���.�[�q��_z��O�G�=]AFHκ�H	C��צ(b��'r�f�1$y�2��@����Y���s��()5f�u��;��$�)��'!��M".�#�%w��l��r�R*��#�/��"�#p�8YjDr,q��a+���m䈺6��i#6t�ݺ[� i�`zz��u.Is��ݜ�}<��]}�I!�����ą�]�
��~�]�ԛA���MA�Fa'C�㯨���}���u �\��6����� `��@�Ӛ]Ʀ
vH�A����&�J�C��i��U�O�@^y=�G*b^U�ֆ�	�@ \W��t��<���L�H�o[ٟ�*��Cv�['<���K�p�j%�;�-|��Vk1�(�}�_�����
��7lJ&3�p[~m/�6(�&���&���g�c�r@�[�u*њ�y�v����ls{�>^�z۵��J���L%�57,	�!���OΦ��k�	�χ�2ܕT����@:280Z�lI<d���F�&jlu�{��B,�Jrn�Ve�:��l�IP=ـ��a�yֿ{�A����Y_uv"�(�[e�rj�p.Kn��lN~w���̨�]���!����c��&&�.���`p/}�
�&��L�1�30�O�G��`�"P�<j����9� ���eaF�LgyX<+�WN�[�raGϼ
����3�;K�����舞��v�4�D�����uG���b
<���: t�\4�(ր2�ڶ�X�9~����BS�q*�0�f��.R��pA��v���о
�/l��8��A�_s�K�J)ʱscԯH��k�����O�73a7�6��U�U��X��⹮&�ỲN!�:Yg7����=r���c	��ۗ� ��E�l�Ud�a���Wk���a� 3�1���g��&D��X~�χ8;�q�k�w��n�8꾲'�h�FJK���ǀ��
4Y�&?�|�ȧ.������2Dڷ�y,y���}U����f�at6,��ʏ�$��0Z��j���݇_�|Χ����N����w���]�y�ԝ���-a�O�`"�[�ō�
���ݨ~�5*��L��P��)�`�th���o0��ᆓ�*i2�K�����5�{ܕloʉ,)����x\{��f��zE؊���蹣�����y�0��
J
N h��R���n�M[`�=A^��b+t/0�z�
��y�22�_���HJPT��N`�O��eO���?�I�u�����j���)V�R3w¾��h�T�0�G��$������F"JZk���#wz�m$!>����m߹���?�`y�Y��v�����`h�����S���!�*b�B��-�e�M%Hu&�^Q�/~s�_a�i(��翨py�k�P�#�Y#v�)�}��
���� �0�>OPz�R��3l>����nP~���9^k�FT���i�U'W��N/:��s�H,/?ta�B��J)41��m<%��W�7���A�y��N%mS]mZQ��%X��<����%?V���xԍ��G0�gy��V^����r~h%��6��xuT?G�?po.�Wb���"{��p#�d�O�)�h�,L�8��#2lOyD&o�� Y����8_kd��5��"��m���c�|u��+7z^"��-�E[Fﮂ�*��v�?ʡ{��e� �˼�����
ꙣ�Zß7T~C�H�?4�o}G��W�D��}h�8`�.-� �ש5�XB�@y+22By_�iq7�K��21p�]ĻN�����ü �����x>x��9������q<\c
��^�aN^	us�P"e ��bm|�)�K&��[
U�� ��<9~��3Cފ)��ҀkX������{�Z(˘$`�����?��P�����UUY�ך]�t�7�c�qڌ�yKd����k٤jL[�7<b���=��`���,��&�i��;��b�N%H��L���B���u`���s3��L�K�M�tX���$�ᳺ���OٺTA3 ��`���D��җ:vxY�o�O��j�� �ئKH��-�)�c;y��4���{�jxUv�Hd��\��o�%?d�{e�D{����݉�b��SP�	�#VS�h�e94L)!���a����fL���%5�߆�Uo���@(�]�+ P_P�SG�6��2��C����T�h��Eh����yݺzh�� 	[��=
߰���=pfn��j�M�\��_��h�jW����l��	�wH�L�0�AD+���!q������z�_�;���#��c��uy腼��QOQq������`T���v���T}X�X����H���4�G�n�c�I8���g]�TL�����6�����Y�}m��[�u��n�b��	/^���'Hܹ҅����o�Fu}*	4�O�!v�� C/�����;�c b�4�9���0:n��wW,k?,�F�P��k����M<{i�+�^���4>b7;d{E���!we��n��զ`��2~��p��~ �����!�i��dC��w�I�]��:�60���\+9���HU��-ܾ8R���hK�@��S�>������v(�Z����_H*t&��u��D����O# �'��m���P&x��)�^�j�h^,��$�s_f���\H�?E)c#�ks�Pѹ� �g�=��'R
	�L1+,ۏ÷0 M#f���=�i3�
�_�N*�a�P,+�ҒAP�%@���HW���Y%w�Dk�%1%!�:��ďj�4�����9�i��k�Uݗ"��h���X"�o]�����x(/1���M��4�

��7m���PȐt2?-��ʟ#�����Ơ5�e���Y=�3�3[�^#A�ق��3��S��p\X��x�:�uo��~����#d.���m�l��K~kə�9�>��� ���+�s%���?���ΙR���\Hf��Z���l;�q�-ŹC�Q���(q�:f�-�zf	U]:��x���zNj��u�wlUir���'D����bG��r��QG�^C�p>��j��]UX:K��BJn�Zגdߌ�Ϭ�O\ۄ#�l��DiH�3X���ʇ���7i�c����C���H-+�:����VH$Ff�;��n��g���*�p��vAiyy�Ϡ�C�W�?�N����$��»����}ef𭸌�@�-#���S�`��Т����d��o�.��.� �	��Y����}��ޝX�htbd�bR�"z�
Ҕ/L��j~��ޡ3�D(�h���A�N��[�����B�dQ-�\{�axo���`p��I�s�I����B�Y�W;y'��_Ę��L��@@Q/i��3Q�GpX/JI_�>���+��*��R����5,��4*������6�y�'�>AB2XT��sT�ߖmt(�0���m���<���$��2������k�۰��%]���1 7Aͤ�͗�9q�@�Oݿ{S�z���������F�o�<�bƍ�"�BT�5��b��O�
���a�����;�������O�,�?�m"Lg1j	%�+j�,�U�g��4��6RU��i���$�� (z��B��A1Oo
'`��n)���|�
�
$Q��i"�Eo:8��x�WP"�5���r�EF-�4���^�{��4P��X5f�`��F�3hT�L����He?��u��y.H�jx�F�̯q@��Ǚ��t�gs��AE`�)�1%��A,ck*�+F_��K`�d��m��e|�Fa��*�����x�b�"/�����-M�H9S�as[pk�d��]�t�\� �4yB>�XA����yw�7��%JAȫ���0}��^25����R�ų�+�k��/`H�Ϭ:��7_��0�}�j�IJ��R��(����_������I1�k�a_,�ۜ��!7���Ԓ�Oٽ7t��M
�@�T"�$!�J�`N([6��7yQ�g`����y��y�|WH�
w�DU�����7,�-u:&ۜ�?��$���3w}%A�$��;�� S�ۜgh!��F'j��)���I�Wh�;8L6��C���� n��J�'I۝� ����ViSڷ�W�@C<$!���Ѽ*����N�	n�%��B"����A��q������s����4���P����'�4a���s��NQ����������v��&���+i	� aG�H<�W�kM5,��_m߾#��8�rW����Do1@U�*ؿy�	+�������7�t�M#6���a�	��BI՚�L�G���>��`r���#�ˣ��Be�qw��Td�|�w��hŢy�<��˭e���JWH@c��|���N��y`�4ծ��hD�I��11�M���&8~�[z�*��e�
�tB�e�85�[-Sӑð�Ie=����iq�>1�uD��7n`��5�.7�2,C�侷9g{�#�O��/O�s�΃X0ۂ��]E�昃V��gl�f��{�����Q�'!(@���u<��^W)Tf�!3I$֎e�
.���^ZH�8.��A!��^So��
N�b4�@��1X� � ����iG�[��w�#�J��.��Di!��Ix���Q�$Y)�.�4�X�`I�*��FD3Bf�]�q�ey�3�x��
��/U �e<kX��Z�Dv�FIv~�K��V�1^���}��u�,/��j���,Xj{Y��g���d�"i��8���f��߮����YW�¸Cd� ��I��I;܉���UK2Յd��$�&d�s�A�ފʯ�{���}o0́�_TZ��ӿ!Wuqk^[�z�mElS����EH�g�;�����-·&�k�ܝ�d>��j	�c,|���ҽ^�������)�l�m�ͺO���V��R>�OZ�j�I=G�u]c�]�1m^�{�����eX���1(�g����c%����0Iyfz���;ҋzI�ֲ=ҵsu(LņH%�����|�KU�p��5���Xy3�f�*H��W"U��G�;�u��>8�@ʑ=�#�3�!�VK��Z66��ތW����20����i� 5��b�d����3]L��q>���Y�Vж��I&rZ��׵�6c��J�3����!�����_�T$��:wM�R?��2r��)���V�SI�̮�f�գ�{4+�?`V��8[~�cmE��mD[*_����\_n��ޙ�u���{�N,[�m� �i��������jr@� ����3�V/u�F1���g��ω��6�a wE� �����Ag���g/�B��-:e���p��2��H0c�DS욇�X��e����5�'{%P>CTQh�S1��S6ZN1�~�_4V���ფB��N�����il����,��؂C�{x�ԁk��Bj�P��O�+�p�;?^��H���y�&6{8 �Wc�!�J�Qw����ϥ��ƻ���@�����H����tz�b���{�%%ݢU�u�~�X�z�Z�6Q괩]8��RO�FM�D6L���f��-��:�ɚ�~^��܋I���#�j��U�}��d��`\�n	naM.#���\�:*B��ŧiz� ��*����IP�Ɗ���-�?=��~〸����q�?M�v��.bf%hv`.��24t�{���dq)_��{�v�x�B�0�L*O�I\S�����7TG.��LB�r׋�k��a�MX���C�Q;����i�U����p��i�i?�b��8�����3���*��>�jo��
U \�c&���z���=�dE#���벁�-�� �Yl�b5BNĲ!&���R�d��U��^?NE7��`rz"J�'Ygu�W����%�4���F�GB`��UKɓ߉�<��}t���&��#�|U�{��0�S'�ܸ����F�����H���reTT�){g�P4,L��3u�d�!Ɨ��cϝ�b�		*��1��?�,SUO2��P��?����Zj�:˪@@�;8o�W;Io����K������D�9��TF�(�f�0�7�]��NA�_�&"!��٭t4=l�5����=4�_��U�P�u�m��Y��F� ۝���9�Z��o5�Y���XEy���e�s�<U��p���|"���vv1ʌ���&h�r�R�QG&��Z�/�����Q`�K��x��	*^J���Kn�U� uC����z��FI� S��o��0GeTđ.g-Mp9�X�]\6CaZ'S�ۮ����?���㕯j��H���Sd�]��ӊ�~���p��fi�W;P�����K�P�R+恲�������3SF����D��
JǕ�
@�^o��}�;D��n�7���h~����ݟ���i�a�u�ζ5㓰�p1�:�-}�8����N�h5�o��N�"E�x�UW�M�c!%f;��ei�t>8]l�������ǧ������Q6�^�K�ve��� *q�T�vL�_��BJ�K��:%
�VT��@��k��	���U�$��%����(.��O����1{�o.�E��0D��xe2j[6�g�I�)��78I���o�oB�"�c�r_֊��PK���p�5�}]0��?j� 9�.O�m-@�.��E��+]&Cf[+���W� �]�#�N����}�<�&Et�s�g�]� �;4`S���q�b��Jސ(� OݜHFp�R8��-JHfɗHj�+!�߻�O�0��}�	?����v����r��l�37QQ->	��n�W��0`<�0�@�+�����CeE�QZ/Y�I�R1�,v�q�`.^��}�����E�By�[��;�V�m{J�)3ma��*2*)���_^�?:������������(�����C�WE�w�	޺��V�2=�]���8��G^��	�|�^� ܘ�#��8!�j��S7�����, ��Bwi�-����š�dr�Vw�Ýv�Pr���.D��.P�p�f;xL,pܬ���!L��a�=�D�MEa�?���9���WiP����k��L����j���o�yq�,K��H��C4r�&S�e7�*��@����	�g�	-���J�s�`  ���*f�[he����'f��: S��2٪��3�W?s�a*�#�k��]��z� ���n��a�Ѽ�oHl���[�j���Ø�V�b0�Sv���2�	��q��g}�J��A��[�EZ���f,Pjt����#�b^2j�3c#*��<(�j�_͚f�e#{�L,�J#l�xO�ݽ9Y\����[�$+���B?���Q3��G��/H��~���C�� ��+RqѨ��KMd�����4�f8os����?)�Q��{��{y4v�Ri]՛�'`��?���^���Ɏ-����"��ϵ���Ȗ�T��k�BD}y	��Ivf���S�(dd.�pz���2��XT��T1��Ǭ��B�6>7��d��H#V�����0�
�-���w��Y��e�������9�q;ո�/��Q}��9jAL� #mA ;D�8t�JXƉyɝ�P搡}5�`[��"Y8��E�����00Nf�Pe���3ʣ���X�`Z�[1-���_\kE�cj��I�0�l�nX-g]ۮ� ~����yQ�-r�φ�>�0!t��~���XK���!I �ow~'H^.�L��~9(ƺ`��o�8{CZ���-x?���ɗ���4��{0�7��)�|��䨂V��Ů��h#�t�Yte�:	%���@�����y�� <�)rv�8n~�Z����X������T+�-����M�����{
"��Ҟ��$К��ZD�  �X]c[�Z�0k�C��&'� �!M�{s9���l^�� ��s���z����0��ΧD���z�On�b�������}�ƍJ���W�d�����԰����b�H�V��S�"͔b��.��A��ܷno3$}ub3�2K�_��gk����Ǻ�ە@�<sT�Dn7�9Al���vw�T|�b�!:Gц�s��,�u�H����j��WI%N�%��9ꄹ����%��mDme܌���ATw�{�LI{ȩy�0y�g������8���9�0�ؽ��6�U#[�9�!,�kM(�J��e(?���R�[r!��s$8�`�}��m�V��(1o]�*N�M���eL��[��!H[�"`��<E� �f���L��5¥�)BJ̞�p��#��,8ll��Wd�#�4E]���׃�ub��T�W��Ѯ/��@7h �M�jַ�xV5۵x0�9[���
����<Ƞ� {l�qe������wǆ)��6Ĳgiw�
N	����:��x����O���q�3�G�|[#Hh��`��Z��d��ٍ�l�5�F�/�0_1 �����oV%S��I�M*T\���ܯ�Y�<�����22+�'�oT��)ֱ�`Q��?�E���Lѳ��feX�㝲�౹f� ���s��u2g�;��9��ϦsT �m�{�4��7E7�+?������R�H�#d(��������7h��H-��h���١L��mF[l()�+�O��J�떂m��0��oz�}��t��*̏�K!M��L-�t̕Cw�|��Du�ۑ���mըJ$g�6��;۾5k�G;Y
1r<nJ�Bd���:�i���F�)C��Ĩq����>���d��DC={�@���\���e��f�i����BI)�������Kj�#�c�m�H��!�!#wU�l��n#��i�b�M��/��}��CQ�F��O�PK�֫�;��-J~(E���=Q_ 㓎6�^_�_�_�b�X\��l���[������v�G��,���m�������t��# �! ޏ-�'��7�,3 ��TP��r���EE���e�B a��"F�����l�L���:�@�-��ôa۳2�uqk!1����F�af���Zlk\� �]h�!��[���pXbe|�d���ͫ���L�N���u�WRǒ���c t��F�de��.ҙ�&�1���>�m
�>}E�Ȏ�����۔>�B��*{)��%��}����ߋ��7?`_�O�wu�`��X�(��l�y�6y��R9}�SYy��wu�c��d�$]�ql�d�)V ���Ag��r����v�n����-a7_��
}s;��:�Wt�ݞ%��
����N���)k��ovR�M]��ZNR���R�)ƿ�a���|p�N���������_�	���>�׼eo�g(:�a��I4��t-��E���&��cd�y~����-�I��t3��/Y�������a~�ɕJVAP5h|մncC(� )�`ɝ�koS�Z�C'ܑ+%g4�ߥ61��ь�rt�B�����d�]@�,O��]y���[d�Q�6;�e��������B�Q�i�%�u�[�:j�d4ekT��گ����X���T����^�M�`B%X U�-Lq(d{a�8�xI���ч�(B���I��葏̞+
�FK{~+0���n����w�C���F��8|�v��󮂚EQPL�:+Տ1�%�y��C���.^e��-����`���
ٵ#K��7v\͘(�?�x�*�g���ŉ��O
ۧ+��ت��ѝ!��jmXn�<�y��V���R7�v>}�{��w�=�F���m��'��V ڥ�8�U�oOzk/g���.���BQj�D��ጷ#Vٽ���`s������4	�&^yVd'�t�(��!��~&_Qۏ:S�p�Fj��25�98L�fLa�d~�r� ^�3���FӁ���#��Ͷ���f����E����l��%k1�(��;4h��|�����3�ƣ�(�<T<g��O�z�1Zo�Wl��bIqB穦�IXs<�4��޴.kr�
/2�S�V����dq�a,� |+�{/�h85u�6*(+l�v���U����b��B�=��q��Xe�]��5�q�*���O>��d2��kj���9vo7�*�B�?������ۗ��/�`�����T��*���X�y=\��_��F�����9O3hxTh惓�R�`wQ�_��7��uA����{$��^6z��`,���X��6�&�S���@c��s)�)C�|a����A�V^˵�O!�)����	���j�&+lƿ��2F4I^,%f�0X��ډ���� �6��K;���/Z̧\[���_������%��ā�_�^�AMP��I�0�Ƿ�r���¹�f~��i='5WzQ�m�������,���r
؄�xa_Ge��R�㸟W0�2���a�ǈ`A�n���,f���Hk��J@Uk[�>M�M�+�yʉq����O�R��D꺛�>a���;Zh�ߵ�,�����Ot�Lc�@*q�y@��2�ܘ����'��ש8�ƥ�C�}��@�[�8�V��O�8��W�����{h2I�|52��dg�84#C�nh �r��9�Tt!�v��t)�DA��~!�1��4S�^�h_����]�cϡ«X9}_�:Y������g�A�G�yO~R�;�j���8ZѦp7����0�A�# )�G��0��]<Zs�bC��c8Ce�	OTQ�:$��WNr���XHZ�\B�S )���<q����*6���-X��3�8�>^�Y-�A,*Y���U���N x�i���h�<Nn�1���_�9r虛���G谏��qQ�Tn"��4(l�S)��M�Q��FT
�>�3B8�k�[˟dOq�f-�Q�LB�[���Ql̘s\k�r!���fb�E"2�_T��ݠԡ=�	���}N�L#�]�����%���~��Ab�w��iц��:yɶ��7�3�Iy@���,�_?N�o�_����9��w�$���.�1��O�Չ�X��W��č��%�(�����8�Fզ2�_�����$�
������{���ܙa��Y�w�/��o�*�ê=���݀ڔ��I@l�J���"B�b�>@F	&�>Œ���O_#�/��)�G��J���ep9-_>��J?���nxO�:��/-��G���&��@�������_$��~1�jG���Pږ�͊���Dj��x+�t�_�t�qs+�L����r�&�5J���Wէ�^�l�����Wvu�9��*ơ�����iGx�' (R7ȗJ���򧓍�ϧ�EFw7����A�ݭ=�5���(���\�ʲn�}ݤgB\�}�)ƨG���d��¢�+o�L�s>I[�uky�h�/��Q��{�`vS#A�L���JV�ʱ��m2p�Hw�����ڲ���QQ����l<�nŷ?6*��c,U�}�gȂ�q��"D�o��V��zC�z��:��<�ʐK�k9��������t�~I%f�j��c++�0�wވ��c0t8����d�s�a��,�����1a��1��_�f�������~x�Nƭ·'"��ߔ��V?��]��re��ĵ{��� g����$ ��ןI���ǦN�yE޸ϣ�:�.�����FO��c�k��y��A$UA���3�Ɯ)��0��R�Of�Dv��)s���$^��Hp����Dt�Ey����"3� z�˸_��_�ȓ���9Cqf�A����R���~f>�9��W�gk�y챮nΤ龖�\�l�r%]+Lk�X�W-�5��v���k��F���.L��c�;=����2| }�"
����mc��$q.���n��^��$B��iB����ЖN��A��ː�z�a���(j��j�LD^wa���?�Qfk�a��:I�4�	�l��R��j�Ci^�#�P���'Ty��=�.;X7\��`q��I��5|���ǚ%X��DT�D-C�hLb�%(�;]�{P����8q�Ҩ_Kp���y���Q���&Ot��:W*4Xr��+Ҧ`K�ٸ�	���!��\��B!v$�~1�H�s�b�8b/z��4���Ƹ x��ۗ�-#tC?c��}�G##t���i�Ë��hWמ14cA�#S��;9�|.��2}�i+��f�}hS�O>釴�w}OL[�RL-���2Ku�r͇���)_��m<���EsK��CP�F���.��t�>S�ġ��b�Ǖ��c�o	���)%�	��-�~j��Ċ��JО��ҵ���	��o�@C�_t	ͺ�&�O�ۋ��npҏ���d��O��,m�~	�)r�-]�R��^���'T�@����	1���(�.���Y ��7X��zh`��!V��V����g����h���W+59��<��y2SJ�\@��wc,<=&���L�_��=�	����;g2a��&��ʫd+�I՚ֻ��.O��㎤�^_���8�+��*m��W(�I���m��
ph��ў/�'Cs�}��.����)@i�C�tT��E_�>r�98��E�������K�D<��%،�:>i6<Mg�������_�@Qr/?<�w��(�,Ɖ���5ik5���#r�DX�3����W��R�)DR�����V"|�%[�m�:G�����I0�iu�y�S�}QM�QZ�;gk��ϻ��W�}I����(?z��F]5fNF��(g�x�߃��S��v=�އ���⠨�e�uc�p�S0Rc���͆�"�J�U ߰kQ�P�ÿ`4mY�<V;�,c s�U���\�Dq~�Kq��9�ͻ����M����ZqVZD�/�\�O���`U�Z.��r^�܎z�6״�r&�s�T�T`��Ik��[Ao������|��p���`�k�}��_��ڹ��u�[�vZ'{���6�Âg���E�<=�n�^u&�p������LG.�7�i������P˫'��R�r ��mŴ�{G���;��$ů<�Es[�a��o���it
�պdm%n��zs?]~�5�<m=� �e�D\ɐ�Dh.|pEJ�$��ؒ��1�DAC����%Y?���ߐ���5�!�$�?V+\��_�
� :�+AdXZӞݕ4 JYc��+����&��}�@
�����0bk�N���1�a�8��"��E��55�=�>8�I�  *� wc �����Vt���_�^���@�^�5`�~�D#�P��ǭ��=��c��x}��Y�m���UJ��B���#7dxt�!Z �ǚG9��F��D��U�o�ҡ�E$f�L��\M�j�;���8l�c��H�۳�h5��=��Ğ00�.V�iӐi?��=��^�0]���T,�,N��-���{���~�I�l�. [k��q@=�(:G/����� �pi�F@�|�n�~�)��a*�|�Ӹf��j�q]���-����K/����WqI-shO�ᝲ��B�z�e�����=rJS���P~BT�'�$��O�q�^+���'�~�����>��!��C��-P��FSrj��$���{��*���u�9qҿ��{���ђv�~�r�$������Ǝ����4$r��P3+�c�r2�~�[�qUx�y.���0ð8���ƺ�=���I;,�y8_�T~��/�3O�#�6�G�|'!N�����9w��q���3��:Ե���\Q�'�I�_��Fjs��ꎦ���ڶ��.�`��4���u�ٜ�Trl?w�����0����Y��b��c��@�?�R�H����X�?,P��+�b�>�p��LL�$J�%/�(.Q���9JyM��`�]Sh�:���I7��b�;ԸiT8U�g�2��[2�hpH��!��MKg�Q������+��l�(Ћ���ɽ�vo3dq;��]����E}�73S�,�!��}:����c�~!�D���E��]~3�������M���\���;s�;a/;y.�C��4:ٖ�,C��t���H�:�?�S�<b�awd\oz"�6�W&�#��$$xJ�#c�k+C:��[���P��'�y��Ȫ��"�jxp�*�p�w	}���=y����y�Y?��s����+¼���tb]"���w�13�m!���]�C�y�}��~�\ڥ�+6Ut��[���Fs �@>�C�WEhX�k�Vl�f1��o������}��#T[,|����Q+�՝
��6I��N������=�3�G���^�׵C���ԎX
E�o\N������J?�Q�U�)��������T�F�K�K �ѐ���"� Ӻ���ʪ3K&��D\���\�����ڣ˟s�zO��k��O�C,�:�M۽�c���Zڊ��_y �.R;���f��B�YM�6@�T%��(���@��]n����,��P&$&)�~j�^�����ӛ�G����h�h�ec��C���i�rM�Qq8o�LM�������fv}�(f�ATv�-oB�Ȁp�
z�*���@,��8�&X�m�7P>��NF��1���A�D8D���f=A�tp�\������Z> E��?�N�?��	e��B4,�L��] �p�H[W�3��E���B��1�؞C��u����i����Tx<�<��|͛؄a;��2�茀]?v�v�Ljґqd����'!v�4`g�����^F��SQ��
��+�rG{N����ǧpN��i�T��iߏ�Q{߂�b�8u(V.ﺹ0�����f�"&��Y��9<}�O<P��\��C�<�����ɦ�6��3����^�b�J?����]��쫱g�E���ir���FU/�+��5i��K6O�ݘ$��� nl��3��f�<c:׺���A��+�����@>W(WZ-��f�ҒoY�����??���Eo�����˒�Sh%xx����|��ZϿE*�&k�f����F��n�X��Z�Zd��̄��CP��j��#���=��y`R�l����#bb�G<�k|�gU"Ju|܈15�uUsӛ>b�S�I��aL0r�%~A�v�QƲ���eryi�İ�9�x��dӅ2�;<:����ȣ�Q��*}���t�_���-���+9u��|-��N�3�z��p9��zv.�!;���2��X�L�!�Ͽ�����<�Y��Yv)�䛨�`�ɉ���+������2�?W2s�&QY�=ҙsde q��} <�}�����T<�S�Rexi�Z"#��'of�^1b��7��%=^� ��Q����OߓP\PH�암 p0�M�38��o�����۟�Ҋ�����v.�E��RJ�9�f����#}|�͐�k�t���O_ʉ��}�'���V�
���zar���w����u$�89g\K�8p}��I�UJV�37m=L01ڧ-"��g��F��Z��f��s�n��U�������n����"-ھ��LA�ܧ~����)t��>�޲|j�ű`��G�Q1h�"�����y��gjԏc�U��� )�Wɑ����W��+24>M�f��vߦ�|��ˮ@.�56O`(��Y���b~�
�<!�h�}�ӳ��⌯3!-�v����I���/r��C/ d3�}-�D%?-��Ĝ��6��׭���,2�`�<��:��m.�&�|+��â����>h+�³�{�0D�o�/:EE�,
G4kD[�X�	��{�q������s�3�UA�g�6@c.N��}���f�;��d��� �}��}���[2A�H�������4�#x��=e�iN�FH�W��}�������ƽ�᠋[�n��\AC�DL2��I�H��xMo{��X��'v?mzb�#�}�%���QYXЁf�B�Kk��}`9��ݦ[-`�'���r*������rr�ċ`��}5$�n�^�/�Yf+�t����ST�ڛ��U�b�
e��I�=���	-���k�>JiA��qr\뜶��H��`��}��Z��V��F�2����Y����y�W[���YR��E1v�%���u�q"�w�k��g�F?�� �������H���,�$Ee�D��	�C�+�/lQ�`j�~v�h<b�i��QA���Ȏ\5��kQ&93��lIe�.4N����f�Ѻ����X0KR7��R\[�xn�g���g�P~ڊ*��̦�@Hg8k�ⴓ4�B�JЉ�ͣ��Ea��ߍ�/>֠f��2si���ts�A�Jw;}����	�K݈Ln��q��D#x��r|z���,%cY֑ :<fcoo��B���;���������=�?
�K;6���֐{�> �B�\�g	��փm.oĢל��)?��'V�+ȊT�n��a�N�b�B�e�9r"ۆ�6pM�a��#��/thL�mc?���ީ,������rg���k��!��줶u�as��zv! \ 5�0�Ы��]k��k�/��T
�¢a�dב5	q�?�-�c�R�D2$�)\4ӄ ���_	��ǀ^��`��U���sW��g���.�p�6p�D��y�f�${��aS4e��&�ʎj��>m�df`��M�O��aA)��T*e�;W:�m�3����$���2�ov@Af��ݷ-��G����\>N���6���T��Pdbb��_����?���~g�:����=���A���Ê�_Tv2�p��2/e��2�����A�:����.e����w�������w=��*}�ȃL��
ֻtL"�iI�-�@��rhP��v����_0J�_]3q?������9/�٤���R�Xt���!o X��������W:������SV�n7�񓧭O���C�� 	�ɹ~�V5����!G=�q]�{�������s엳F8���`�uXlv\pn<�x��_0���dAY���l4�	��@��g�6�"���@�[�83�P���9c�9��i�;jYF�k
��Yv����U�Oh�ε �sC�|L���gƗ�����8%O�H4I�5#hyd��ݽ�s��m��ˑ۴�WZZ�dHf�E^�d�F�O�Ϲ���o5Ո�"8�W�l�4�J�2 .7���S>!p�?cSn�!vQ��H2�?�/h��8�w�����x୮t���&t1�3�s
Jj+�}?:��
=,p$���y�r��v{A�Be��-q��2��Izq7]ŉ�R�قςp��`�p3�F&MT�6���}���jᘢ5�S�(�-9�4g�
�t����d�T���ܐEq � �b7K�K���=�q �KV�s�
���e�P�ղ�~�de��ܙ⪷�܎n@:�&x�q��W-OӉ'���@���j�mit���<�Y)x	�sL<ԋ�y��"�&C�]BǤ����T܉�f{�O?J8��b�:�Nu
�k�Cɇ~�@�̇��F���b���kt��v��,��`stA�$�k�z~�tS-���5~�!�u%��zNܮׂ��Jzؤ�0PG�l���&n& �x�������Vݹ[J�خQ~�=k�A��������7k�4-�e�)`׷���<3`����x�s~�_��p��cl�Ca��!��>֟A��I�bXこH����i�%aݟ�獟�?�NsD3Uҧ��hP�m2Q��<J�&�r`',��^ӣ����f��a*Gu�R��=*� -\?V�V���՞ʀ.��b_�G%dF������K��\��Q� ��7�^$�����Vhө��������Ӂ��(c���SG]DٍT��yD��;x�澭,I�/�]�8�T�?��Ց�N�� Ň3�Ur�#�m��Oc��e���EVIͱ<��l�rc���q�{"�%����g��2���X:}HqGi�kM/��عf�)�g��V����.���� n��cBel���IN�l��-��d�l%��� �nBkh���^���	Z<h�1�,�DS?|<cf�����x�)��!N0|���s
���Fc�Ѭ���D�Ƹ͔�tD����`���X���noz�V�w�&F#e�_���bJx����A~<�Ö�m)Qyj���M���/-��
�=h�+�m�CǽS^��`��N��a���TC쥐'�A��	�����G��Z,n�6_h�8���/C�Ր��g�o�}ҟ�m�;����t�0V��lw��`�7W ˋ+�*�}���R��]0h=��p;�'�poO>p��?�����J^�z��~��u�FO�z£�����{��>M�4O���k5�cQ�irj��k���P�T���;�;�7�,5����CQ�{�B���	��aA�Z��
)�"����iʔik��L���*�,��K�6���k�J�փ�-�����^�/����*pl�`�KzN��E8�t-���}����E���#�Vw����f�{�ۚ�0#z���̪���r�:�L�����#2�Ɲ��y����u}ĵ����mY�s�Q�>%wb��a���#���)�޻>�W�N��X��ǱP�x�����XCF�uj�P�x=�<[;(��t"��?M>I�.�єM���.:�H��}�h���S9��v��,H��a�
t��1sf��ҳ�"MNo����\�U S�
S��CdtX.��QB�uV�%E��Od�Dp�G&)���>����O�g3�4 �}�S@��d�%�oQ��#j�Z��WB� ����m\�_$7�r�6����*��I����N17S���pE@j����ʱH�|�b�f�`�T�n'8Ϣj0*��i:��ʒ�VЋ������#2/�Ȏ��9���:�X(ld�`�������-$��^f��7Ƕ��a"�]A2� �J�J�W8���]���)ԕ������-AQ"+|��OK����v����}��AT��ֺL=�a�A����aW�D���0�{���(�;L�<V����ez����b޽�Re{���^ȫ��W&p����lڬ��W�d*��Y�pL�%;U	[s:kdI����j\�Er�ɀ���WK��$@�{�O<o����c}Pb痫%���w�ǧp*9����9��#�f�S�F# ��w��fװc���Q<0wmԪ�<��_�����P��e�xL��@��\�D&�g9}u����N�OBC[�0�wٓZ{0%��zd��dc�j�h���Kc4 ��}�u(dH�	5>���F�^����V�n���Y�b��x�n���6D:��}I�I�6]�㓺���ɺN���W1�./}> ��s</2���Z�+o���=�6{�X��-6"�F�2��W�b#�I�Mv�
���C�t���
\�}'�o
%I�k4�E�l+�mg8t�l	�����m���:/�_E���P�5-5~v	۽N(�K�d��ǎ)\GQ"9�l��R�! ��L�����h�HŻ�)&���������A������T �eŲ/��l�z<*����Tm��}�����T�$:=9�����Z�ТT�U�~wǜс}۫"���MS�{Բ geT��_rn9cM�.ɸ ��/F( *)�ݦ���xl�sJ�����pˌڥ��ᓣx9�*�	����S|ܫ��~�>�;��!en���!XMZX�^$ء�3-�af��0yeS�j�� �� ��l�FV���;�=
��.��U*$�W<;|�Y�k@Q�a�vK�o��sBu��vC�|�ѻ�U^�FCɣ��5���ԩl��skpl�Y����b`�@�h���^ֹ������B�#�8T�}��e�V{�kv=LEjku���޹��Z�ik�l��1��~�L X"K�C�ΖS�;�J��Q��8�~#&�������n�5π�p�X��0�'�q{�4�/�Jb�4+]�;l��`ݏ��Vĭ�H
��]���W6O�����ŃF�x�K5h��o!�֍��*�GX�Ю��`�2~s�^���X��[��m�#�Q�:n���
�Z����7db�.
��'���R��g��(n�S�����%L-S�ʾ�4���q�s�ҵb�[S�)�e�r�w��i��贆^<(���{��ä����^�h���$HC��`�]r ����%	jPa�H��@3�
���-��O�+~��gi�Zx+9���0i�5Xo����{3��@8t[�\������O)�t�d�ȳ���z?LZ�5�/!�>��)�ɷ����[LY��Ѐ�ɺgp��m��;O^pu���m ��޻�S���p9�a@�:f��>���rYXR���&6����z�f���գ�g���}d5 ��+z|$��E[���m�?6�6H�֢��Q)�P]���A�B�����g�8~H7����?�n"�Ƈ�~�S	d����V�h��r�3&�Oy���~��h���V#`���7��v �^���`�6R�K��w��@��Sʯ��KI�C��G]���Y�@����|�Y~p�K���`O\h�_ؒ�m�~��5q��$�H�G�}
��ʞ\�'��'4V��u'(�E�<aq"hg�C�D ����w.��m/@M�Vj	F?4֟h.���d��<1A�R�ir����f�n���z�C�c{�G��% 2�f����pך?i�c����,^j00VƖ��b&,!9b�"5���A_�G�Rx {EG�n���&y�z�D��%*�g�wz0h�����I�qy����g�z	p2�y�8"3ш�,�Z*~�YK}O/��}-�IM��
>�a��ZIj�k�>,|ϟE�6N^2Tn.Bp��wL�6@�tb��U��T�S𬀭�B�A���M�������ͯ=s���!9�0_�����O�i{[vb怊'�u� ��l>�ȫ��D^����m*����`���:?�f��~Ozq\T�� �%Y�m�����ƻ5��������HmB5P���d��9pW"}�&Lw��m�J��"ǵ҉�l�T��܏d��9Q�U�B�D��&�����k�wbt�
� �\�{9�5yb)$:	F�����h
�6]�����M�� �����V4�
A�� ����b �6������E���/0L=�D��l_!����>����:��Fm���aÖ#Kk�����P�$�
;Cr&
����J$BS%`����6�^l]��5��:۲��d���,�d��Z"Uc7@'��Y9���3T6=�wQH���[�s������+�7(��p��	����̊���%O�^zL e�g&�"NG ���󞇻b�bQǂ����;�c�B�<C�l�������l���~��=�ו���Y���m�>?��y���qr [a�Z���4caC�ێyǛN
(߭7�_-d���[�qbƲ,�����r����-����<�-�P�Q�G��~%����7k�i�5�x ������N3��i�j�� 힞�LeP��l<RUT��r\f���xeѰGmt�fӴ��V�<��N�!����I��s*z����.�IO1u	&?}-an�r4�VYF!rP��~DT��=�unҫ={䒭��g���Y:�dT�;v;�UA�j�%�K<ώ��=�6�Ǟ/O�\I F2� )#5yc�.Qb��/0$[�4�π��B*�>����`������%	��/�g5 �>l���9��G]�9ڲ��]�8.��U{K��'��)�WO�?4>�0D�γ9��e�;�H��~:�L'CQ1VBАF�r�� �#mR��Y���D/
�4�M)��Ǌ���<AwhE�y>�{��2��B!���ˢ���)c(�3�O�C;���ɔ1���|�{=pz��qRN�L�)[R�نa�N�q��t�{���*�kg����EJ�.l���Vu�|w�zw@�Q���1��\�����si��Ζ�\�At�~����I��z�R�.� k��J�y�3+ ��20fG��� ��Q)+E����h4C+�P��ѡ�n��p�&���M2֌�CY������e�_͉��5�dz��c�CҮM+/�
��A�K�NMy�x������H���8g�A�-�]a���ٱ��F{R!�d��4B�7N�Oi����ܥB�9���r��p�m��t�c.-���"؂��*:aG�BZ%���}qT����t�7���e�3gu�Ȼ������T`�w���}sþ��;n�Xu�%�w���q�9�W�؍L�V��`%-4�%P$xX�$O?M��*�<jI`.Mz�i��7y��P���琡ߐ�]�)�c��m�IvD��t�����eR'<��>#��#�t��������@���!=k�~��U7��N�#R@�hBL>˘!1-Q8����2��á'W/���>�1���X���Xw�h8�{Ґ�5�p_2�E�������m��;lߪB��A7��ل���ʬ3�E�r!�N�Y�0گ/l��w��l���� ��c�_B#�T�B!�a�zI�z1�c5L4���1??�M����W�y��y�l�K�����?}����ñ�l��R> \ZM�Ǫ̡z��zn�E�Zo�3P�Fry���)eh	%Jp�
��s,G�ckHz���yC��"-3��y��P����������u�^��I��p�l{D��"k��ev"Dؒ� Qès-?6�>y��$؅~.�ƶz�n�Tp	˽b+� ��;}�n���.�-�t�)�4�G+GC�U)ֲ7���
��<����35x&mw��S��8�jW�T&R�@���a�w�"Nۥ���y�Z2q΋�4 uZ��X�����&�ڏ�(��]�i��6jr�� ���+8c�Y,@�M9�^C�{�Ũ����|�av���E{�|�v�����b���a�p��6*��Eo%BBU��.�Z/r�������(�́:�{Z��W0�x��M/���K�%��b�Eш�޵R��В��o��?��^%�5�$V��̱���0��:�X�,��ʪ47����8�[���i� ��:�P�c/t��o��Bɱ��U��xU}(����ڊ��Uh���ܴ�1��.�oQ�y��yҴE#�+�.ku�_+���?Tz���Ŗ2ԕ�([�6��?&�-+��z ��-a9q!AI�W���+�4�C�>�ؐ�O�:,�+=���D�Y\u�/[R�KSMܶ�?zwk��X�Y'���D��:��S���~��.��� �l����x�b(�+C���+��,��3�YNU�<)=����s#��+�^ ��T;`>1���#X'T���~�����ί=P�!a���K~l[�@wJ?c��T퐹q�t?��@����ޏ�1��`��;�O�@UaHt�h��|�衇~��
�E<���i|�]�ӯ��|�ViI�|!M���X�����Zm��K�����S\,[f���j%����{fmv@��76�p� �8<)�&����<$�_w�[nME�I����ݚ��IKÕ��IF�!
R��t�sX�<N�Z(�P0]���9Ju�P�0˸�k��Ex9����vVl'	RD��>�o���6�!t2hRD�sp�NG~F0,����'@4(��"+�Q�������=�HT��(����bF*B8o�E1�-
��G:����r�,R#r�IK`�.s]�A-�q3�C*����MM�$El�"�2��h�5��z�R6�A�M%�V�h��Kb!D��sI�g���8�uM�1�b��P��jP[e��Pu`�������rP~[�������a΋zs�T�&jA�KѹJ��P~]F��C�x�hk4~��a�!�k:J��H�K b��`0��?���\T��y�L!!��T]!��px<'���aϩ��5�k��&��0�噙��lo�e'~Ba`(&�����ګNՍ5��P�d��잆0.ay z��ٰ�ЇU�;��&*�����ZtP��a�� ~ۧ<íG.�p���|�bɏ���,8�p�?�-1�G�ʳXY���j�Kv�0��Tt��)�4���a� A9U��وJ�����1�O�ws&���U`���U ����#i�*�qİ���r���YȦ��t@�!��:5y>�]3�����C��j�a�D��=J��R~��
Φ8����?��mB��U��-�p?�.q8�}�^���,.M��k&g���1.��=R�ҘOT��B<���f����j=?\�2壖M�l8��d��B�z��<}X*��\/�պP�(gOl�e��wkraE�ׂ�l�C��N�f;l��H�P �]Q�^#���?6���Dz�4���Y��V���¨�P�j�7ڙ���$�B�*�jD�)$O-o�rG��y{f�Nj�L+��_���T'< 7���`�ћ���}�$eF�)��[U��؋�S�|z9�.���6>�
��a�ҵǝ O\qi�L�H`�G!5~|�����͈��/�}�Zr��^秋ƴA�H�a�BzW�z�Q�p<Бy�I��BΗ�Iw�;TN������1Y�O0Zv�P�c����Y�� ~�rُ��e��F}7y��E���+�&��C�	�aw4z��Ca6smUJӚ��R�H6�PYc ,���ʨ[/m�ڎ.A�Aܝ���a��n?a����%D�'C���F$� ��R1��+eۭ����Y8��|��1��U��>sMn��|��m�>�AL�����^�����;F9�l�Y� �z�%�J����b��]�_�wO��|n�}����|lJO����i�6�5���*�:|rѦ'�[=�k�ag���D9G1�Zk��xs�{�)Kz��!��(�xb> ��Z�Wi�:+�ן��8��L^���|ɺRW���'�k~����E�P�97�j������bb[Q<���C��O2ͱ!z���%�A��f�����̙=ѿ v�_1V�N&aך��	�r*�-�U�b�$M�{Z���CR�+�>�M\�i�2t�C�\�:O�G�r��	���󷔥`��k�(~��$e���o&��o�e�N��O�,<>%S4�8l��]Ӌ��� ɳJo�<)T
+	�7���-��#*~�)v~��$,'�E�u��P`�/�+��~5�F�,�~�� -�����h�i�+�jq&V�HP�����Inw���W'�{�H�5��A(\M��"~�j��x_=��]ç�9;��Ǆ=�
����t�oʾ�w`�vM|�~���D��k��Կ�g1�=�1ԑR�}z��Mmi~]����p�H����j~�5�y-�ΐh	�/�D
�aR���N{�~m�u��i�������<��6B�OyN��.^��py�W��y/���7bGhj�߮{�D(M��2��کʣ�z.��l6ə���u/��y�48��U��[�E ��E+y�Ս��a1e�8<���]w�L�0_6�+s-9���s&�w)���cӪ��c�4��o�D3�����'<ȱ���c���-h��"�l�,����Pz)�q(�$��i����������%��l#�Q��!ٞש_�5��ZCO/T�Eq��}G�P�F6�;w���>�EnJ�}a��_�#-Hrq���j{md���iZ�1�����.���8��L`�P�*����V�;�Sn���2���J��PXĝ�f�z�/&����PR�������]��&}�i LwE�������)w�mL�ZU[�v�lȷp�p��j�Wj�	��P;�h��{��&�)hMy��T��y��_���<�M �˫F���T��ݘ����h�I�=td�[��r��
	"�X��~�m�wfeّ S˕��Ց!���t��F��n���"��J�Gj�'��e��^� �d���k����݊���A�YΉJ���;�V��z��M�՗�s+�X;��|4�ܒ#������j��p��W�I���;o\E���z(E�� �xkZ3:v�z`�N��5W/-){�=y7�;�k�UB�Od]!7����p�7
��c��TkH֣�̳���8T11˹YZe�C�*�w��@��6V��0�L��/U~�G�[ʱ<�\gw��Gx�.u�������V��g8����m�Q���}:l�j�x�΋���<��	�c�]s)��:IZG�5���W�Uf�� �}�՞UO�yIw"[w�LR�I��	�i>����Rʫ�Ey�?�3c<�`	G�G���|2L��l�a�qQ&�%u�Ԧ�3��-vO`u�>�{O%c�+4��*�|c�Lj�pǘC�O�= cW�	���BR�+��Ȩ˹�!.9��G��RRWv�!�b֗�q�FXO�X}�/\>�!�I"��KR���S.`�ⱕ@��܌���,r�,m FҺz�?&2�M����e����nB�G�r�H��@D����������6���B�*����n�z(���9/�3�]�����K�����"���%Fz�<�PD����S�8|..p&��?~�F�Lx$1�)�7��Јc;,Q�h	ğ��[d[#g5=�n	���%5�,���[���(ޫW~�'�Lr��^�.l�2�����j=۱%��
���)�X�Eotf�e�1��z�Q�f|�"�	�u"mc�.W X$�!�ު���� ��5G�1�	ɬ�j{gka�o����w�ɇ�c���z"���w�T�6i�́����Z��8]��`MG�&6�eB��4ͳ�#�;�s��7��. w�ǽ�B��Y��
1�|iA�MQ�|��v���Ԃ�s�X �?AC�0;�m&�Y�y�IA�w�,} �h�\Q~pܬ�m�JåU>΍=�b�O��Z���a>��Q1����U���2Z�kV���<G�B�%���g�n�A�+�H)y�Yw&�0R�b��ybfϞ��I�����F�,j0�Z���;��ư�b+h�ȉ
�F� JH����wh14G�MM)A3@_��f�|zP��5�����:��-t-;������w�q�5�׃B�p�e�����#�0���x�����zNH.&��Nv��(����4������{ k��hj6i�~���|�^W7��~
Uj7xkL�$��ù=s�8AB��(���	f���lYWͫ���;�� ������,d+:����vt�����,mW;�_�<�B��4�	9�\���?�I�'t�gO���� �\�D󯡉�$��VyJz_���ͤ�m2�)��K�Bv.}���z>�B�(B���5I�>�ԡ�v�oY8��i�{	́��ߓ&�nL���-��0�&I���]�y�D�<�z(!~�A�m	%����}J8����Bʪ�m�n% �T���������q<h�B��	�R�ZB=:�>�ǵ�{'D
e�>���[�?cI悚����K'�Wձ�`·��MW�]c��sS筵��gq�o�M�y���5mKP��T�w�Ym����Y�ٸč:t:�B�9�de���>�}���{{\�b���Т������@4&�b[ڴ��H��BX���|�B�����Q����y�fe��ԙ����pL��m�WSra��aU��?�xӟ�8o�t%h���?�W�)dEsd�_KA���I��@w���g�Ɖ.�1�Qn��@�J%�M��R�
�'T�S>f�S&�'����)�>���
1�Y�\6lu���Ӧ���Y;����~n� 5� cۃ��xy�~�lX|7�/����i�����%��V�&t�m��zc�@,��݈���=>N�{^�7f�e�;؃�Oe�8*��ʙ
J��a$�p�e�K��� �X�}�SoV\K��_�#PC;��U��jF4A�W3W����0���<�6+X�7��:�w����D�����G�q_�����͍6��j���B��-)<��i���i�T�&1+�`P��H�M@hd�.������c���[aJ��r?��p�_��}nȘ�T���j�t��k�u�@.o i?U86������!W_�Y�sRJ�$|���c:Е"��hk +3::b�_��]��7���h��`9o����\M*�#d.�fSϊ2������/�əA�����K���+D�䒽���o[IYJ����o,���U�Qq�$��=� ���8S�L*q�v���#O����H
R�A8K���-��Q�շ�Xa�_��'����#"~LWG�`�.��x�L�X��;���k�My�.���4����Hu�0n�;��V_=�`�-���m*�fcD�V��Hq��i:�n��6G��'�S^���%�峪<�F̲\��k�
��p4��QZO����~U��L�����j�b�h�m�{0c��N����gA��`Χ������?䴎�
%��}Sz��-/I|��7�L��k��C	)��h%r"�%��&P�hO�q�EFU~�)��9R� ��*��@͑-�+>�S�NESYzLg˄'a���F��m�䓥� ���ē����|��G20A����	,n k��3�S�e��$с�4,?!��s�W:=��Z-��+0�9��MM�8k({���X���XĖ�5������P�$]��Q��HK{�W��c"�=�̿lHz�,���3C��,�]���5�G�Ϋl�>��ѫ��`4@ &ŏ̮�����F���O����z�C�?N�����}�IP7������Р>"%��9��R���d�f��^vl�3g*����9�9�|;��π���FiD�)�ԍO@>�E�����sCXLx����Ӻ�D��A�2x����
K��lM&�A�[�ӂ�|5W�T��i�c��)*@�)�# &�&zp��{x�Z�״�D�?km�ѳE���O:�|��\(��')_)3�,MH%K*�ΛN�sE���k�?�a�?�*���d`8�{l�R&a�w���m�u����e�Y
�k��y�h��48)�r2�H�l���.w�$�:Ueh���m��0�N^�vo���Cv�����1I�� E����H�<�o\"��Q���0�s���EkrI�BEi�d:�&s1���R�
�w&�Yg�qč{�;�����e��}��D��};��b�JӵD�hbtA���I�>B���lR7��A����rJ�_�4
���Xa�#�I/%}�5�OB��m/���c#a/���k܍ה*T��`����$�����J�r��8����\�⎦u<��hyD�+9�o_�A�L�Q�׶��
M��;{A�]'>��3\�]j%qLV�&(]b���|�����$<�)�Q%�K�_�i%�p;�*&h�J�����BXN�⮢�$�ǈYG&��E�	X��;����� ��Ä��D��k㤣_�ϟ�|�f$A�|MaEr|}�kl`�Vi�����r��q��j�h�2{ U�=d3�Y��{�|�`��:G� d�H��G���������h�t��g�*�R�》�|&_�ȖS�?�tvY��� ��J�F�@V�q�ml��a�
t���zysn��W��%/^�c�o��y"���)x� L7T�/g�L�ɉ����u�Q��1���5�\��?���*'�B�I�e�{����s�/#���zC�&1�r��;Tmcjשe80�S�n.q+�����<��:p#�a5$q��W�6
������m���$D��N�Q�^V�F�V����kK��/0Ȗ��
��Lr���~^�ʵh^�9H�^B�R����܄��F6���~�f��w
^�zx�E�����_�R��~;o�����y"�k�ͷ
��i�Y���A�{��`��-m��bi���44��,z_��^ �we�<��㷞8�4� ��XB%gσ�Q��!���_iwF�@��v
��'�9���݉�[�J���S�&���j|���U�y��0��&�t"
��x8{�/�C�2�{��]�)X7Fp/¢j�;��
������n��Rӭ���S�1ݥ�Z���k"7�NUDG�}��J���b����/!`D:���uЕ���6���C7J6�ul��	԰jB�:HQ��s�e�ЊV0<"��+|�Z��ș^ Ұr�:�f޲�a�f�?k0Û$�Ա��M1[�2����P�2����ui�X�՟���u�Q�ƾ��
;�e��`�QƦ�B��i1�� ��_}W�;��V/��=��#t����E^dx���Ys=���;,���׳�,�X7�'_*��r�4��������R����8mI�)EioD\~z����C��;���l�,��cOD)��T�
T$�Z���!�Į7]���ot_Z_)�"����P���.�^R�Ǜ��Z)}.2�/#͘��`���X�_}�
�z�j��'x�c�?/K�jwеIXW?u9�(�� 	�"��G�*�
�R�|��-���b�O���:����k�vV���Xe�"|>��J���,��-�1�&�hc>�;z���rqq�Z2c&vpk�{|����*Hv�-���%�{�%l����,�َ�:�	���2�p���M�Q���q�JjU�=��P�$n��n����5���>V��2�G�	b���E]�vp�*�`V�����λ6��sYZӶ'��t!m'�|�ߞq�oq�&���Β^�d���X��@�'�zq�����
Ϙ����^0΢&]B	n2h��r������U�)6쩤���ii��{�`�v�=(��O�R�n�Á������,_^�����OH͢����TdpJ���\ɉz!v�\�쿊����C{$�g�32�?b��F(|e�W�|Z���l���ﭕ��0��M���I�O���T���R�pr�������ҙLA_L+2�(Ԓq�B|�� �[X� �+�G�Ӊ<��we��Z�1�CyX����8��l�ZX�����`$�޼aҲ ���і|���~a��Q��P9�Θ3yN��;�+U�^7)E�^����⼝P�Ծ���TN�l�qHA�;��skf6�1���`ȍr�#`f-�9��jn5�М�6��l^OX�P�UL�1���߆��Pp�9��#N-�S�F�%3�������҃�^Ъ�q06u����]��l����v�m�y41AiV��Y�K�@���Qo&��v�j)�״��l��V4�
p�A����#���P�n��`�=�}7/.�Al�7�H�f\	��Mb"]�R�K��%hʣ� ��I���V�-��njZ��� �7���&J%#W	��A��`AU�&�vJ�3��4A���P?�峃�6�\d��$6�h�]b(�V�U��m�(��M�6{7kL^O�?�)9���w�]��Ηg�j	ԓ�V-�ԴZ-�H��%�,�*颹��ۊ����`��&�i�'��ǔ3���q:��ګ�y�h���w�J��W0Kw2�7�$��'\,E�!��Y�0��๲X��h��a.hUsw�Fd:�8�#�1͑��lN�u�"5��&�v���i��"T�+i�#��NRMx�34�g����o�Q��I� �������"�;%�T��F���`YS��SB�x����Q��
{��8�v�0��KH4��J#�E��OU�|>�6R�,���O��,��-�0�oBAL���+����S"^�T�	�+�u���������7yJ״]��	�:@�y�,��Y���I9�s{<��_��ā�;1<ztLPM�薩=>���It��YP�dq�Rǣ-��!A�qZ��يIx�hI�螓��J�I��f�#w�ؒ�����T���(TP,jr��7k���p6Y���V>��"��&�P-�>K�$��Ώ���*dt,�/`��NV
]"8@��ھ��s��ۗ6n^OH���W�Eg��뷦�]B��n]Uzcٹo����j%E���� �6/@��U���u��W�u�f|a��ʢ�;l���^���cVs��c�t�������J�X�}�f��k��%�Eb$W���0:�5��n�æ���y�^y@�˵r�;��5�P -LYR{�g�U��1L���y���Q�Т�Y��KL��$f��G���+^�����j�Y�` �\B>p��^Qi�9�����=[Q!�NQ?\i������J���R�N���[��E���u��t)YD�ދ"%t3�	�)Rj4�$T�4]��#GP�@}%�/b�ù��e߹���W�B��'3������/�w|���rr�G^����gws�-8�w���m,QA�y��b�3����?�����uS�C���=-b��q� ����$zJB�Z�GZ"&-F` ��D!�2��5�B����5K��)���(��Dv�[U�E����=�C�)�/l���&#�ZW@1"�@�9�-�~S�vdN�`�3؜B��pƁl'�6��;��/��A�P��:�pd^G�Y��,1��b�����aB��aY�|QOl!�U ���K������f�h��+H���M�8>ȻXT-r������N�E��c�X�*�0�,�,�g��xvV}tA�~�$n�����hb� �l�@u�X�t����O��f��_%v�N�����<�&�F)����~_C3�_k�,�k&���7c�)Jg쒑1����|�r�UH��D�O���y���	L�Tbj�g�5B�I5ϡ3��Ϟk0��5�;F�񟯕��G��U��V)�%��m��;���2g�s�+�A#F~U?���q�����d��<���Dʚ�A��}X��͒��k�)�؇a�C�S�$ʟY�a���AP� q�w��]zf;��$��9�Ru�:B	M9�m��\N�״�aԷB5�����}����%d��.ۭJ2I�z\|*�j}J{���]���D"vcl��|�9bD�Q��ZV��K ����w9P�b��[7	Q`,��4޼�@MV��>�M/�'"��7w�e3����ܻ�#��L�"�רE�wӀ��iJ�r�m�����{\N씒�~�Iɥ�@���=�$	�e���F8�^V�}-c���*	[c�)F�T1�Y�Wd��vl�*.ǐ['ߎ�;O�G.�L9yC�@��$�Ĥ\XOA�嚬Ъ�*��Z�x��a�+�U����yS\'ę�5Ϡ�hB�>��>t�J&�AZ��@q�PGn ݘ���Ĵe(��M=%o*���.|�;ė~n�(�%�Η�����u�t�t���?�5��7�Z2Z�zZ���^2a��Uo�ƒuj��"�p#H��9��F���� �s�g���l�)�G�iˍJg���	�*
qk%7��c�x�t[�`/�9K��0�&?	mq0��R"��^:/�5���y�(��p|q���9�a�~�>ݓ�Z^�h�����.�n9��;Z�����*~E����򇴎C���b�tKb�F�<�+��� ,[k����a�k�ΗR4�[��ܤ}��Ub����8�	R�F��Mۋb�R���G)� ����#.l;�#mH)e�Q[c#��;3f�&��y��N'E����~­������W�;+�b�<��ss6'�@-�;�,S���v4oҳ#u*�_�w����<M�W������	���.����D����3�iڸ,���J�tBU&ӫ"wvQ����
��/Aq���"S��l������y�+$K�wcw%>�G���M�c_��j��Q	k�5S[?���J=��8���ˎW����1w���8��=I����)��>4D�4����a��^�Km{�w �P/��}^�gch�kØ"T�{��ܲ�4������9�I@��c�t�'���@66�q��. W&�N�������(���ꫜ�P�H�9��x�c�-o�z�?wT}���<;1�:/�x+L���*�B�/;����t7s��w'9�r�"ƁQ��������~&0,2��V��6�0I�r4�tw�q�d	D%�
	<ѝ�չa�]I�X��;lSm�����ٙ;���ė��(�f'����wNt*�G�O�:BS����ٕ���a4�g�1F.Y�lURﾅ�ɇ�l$+4�)�4.��E�?_��
�K����O{upO�.բ���
ݭ5~��j�L�~3P���|�͎���J�Q5���[�-3��83�n?}�"
P]�2=V��$�:ǙZx�O2(o�i�D�X�j�C�Uq��~4�u{Ԉ����_w�y0��;1��72EC>���(x�M��d1diX*�)�7e�'��#����GH�F�&��)��f4A$? �bɭ ���#wI�^�"���ĉ(�K2x�=Ťu2"��M&�F��Xj�eob8����Qb���@w-'�o����m�zs�����m.g3�驫�K��{� 	������i��X==7NW�e����W�NȒ�,�C�˛wK�����T%��P]�,ǁ˛�/WM~Nӥ�
����� We���l��{�v�����g�c��eNu�����	2c[�s-��3��uB��.魳';�=:�t+)v^��"dȦ+!��r��F>%h�Y��@B��lNy0�`������!z��Jw��֋�i��l��}|܊��!K��-��`��k�-2U��D����a�h!��@2�LSķ�Ϗݿ ���r�K�ᓉZv(�<k9.��y��s�p�KM[�~t�=1�gl� Ogk���kp���9d��>���L��EԮ�Enp�|쵥�����c��As�C���@MP9UF>��Z�mt1�2���w���iPr ���A�-�� �<z������8����7g�����6�F�S1:é�089�n{�i�����y0�hڷJq�x�;Bl�W��쎜6����߈] �I�}�s�C<�[��:/����@�P,$6�F�x� �hT������Ye�$؇���k�\�=4�t���G�v��N�xe#�8]��6����a��i	���Kz���f~��{��G������K���~���=���-�f��>�c�8�x�7�� �iDu	Wb�l5O,���,�{��L��vo�y����DA�"E�;�Y�Đ�����h�ۏ��=��;�O������B$�s��hm<��7��4z3%��)�Z���ٴ-p-�ǁ��=8�@�$wVZ��ǒy���Jjl	�q�W�V�Fi�lU�jS�\q�.09[K��y��e����^�<���	��S*G���\�`�X��,ͪ^��h�~AY$��R=��f�;���
B��o�˽�}���Bruҳ��]k��P2_|"�q��`�5 �R�f�8�j�6ؑ����=5l�c�~o1�óVP��hyV�9'�n��9�*L��M��%��hBtbzа���.����� j���5m�n�l [�%�/�a�#�ؔ79;�N��!+�����	>zC��J4��.!N����N'�7Rd���O�l�s]G�?����qV��5�֤�V���Vml���F7�Eح�\ِ�g󼕼�~-R��JĚ�^C�@1�(䘂q���?���L'9?@^m���/�*���}T�����N���̛حc����mEֳ̙�vt��p�{���R���ԕ	���� �<P&>nLv���L�2L���I�$�(�_sc�g9�~{��^�G����'ZU�7)�E���ǱE� ��],j��)%�*jo�x������е��_2�}��~M�)�����C�XP1�m�G�[�`�x���o�Q$��V�i̸��ۏ��X/�b�1h�0H���1����g?���06oє�i�����S(dY+�t�����]H%�T1�9s;�G~�O�Ǒ1�H��=��dl�}z=�:m��󤝼 f
=�a��$Wx%��8��B�Yp��[���`��ޢ* YX�(�*�;��ӨЄB���Շ%G��w�m�$Lk_�:P��� ]�+n�T��H6��s0�r�y�2��<Fmr�i�t��4b��F"�}|�gc~��E���Z�Z��?�	)\Hyt���Rn�M`cNB��j}%�J*Ly1�%�������l�No��`��.S��p�	P�Hѓ��d]1�QN�#�L��Zz�����R��`e���ʗh��{��j��
�u�b��m nd3@�ي�Tf��"����'.DW%XX脆�"�Qg��\L|@T`���P!�
�oKJ���\�H����"��"o�ȄDۣ�QQv6.sS0r,E�|`�������vr[2?�6q��q�~h�Ē�2�w9IKw���V�n�ő��+R��*'X&k�����l�a�ż.�� C��N<`_�i�֓(�zI�\}��2�㮘��f��0��YM+-Ԍ�9�IWS�8���(8���� v�2AN2����.��[e0�3����0y�+Lg���1��V�d�tjE�n_HT�d6M��9��e�X)�CͷB�>X��.���h�I��}��֞�e���:�#��9ǲX�8R������(Nt�����-t�5�Q�Uz���� ?@�{k[RyȵF�^��=�F6��v9���C���7�=�'����1����Up+Ծ�s,�ۆa���������[���5ΜG>�G�	�s�<���Y��P��\����u8N�:Q�0����Y�B�N(�J�6����)yO^~������e$f	%R,�+�ʿ�j��_�rԔ�e��OJ%�*歕g�M,��)�`O��2�D�M[�4�5"R�x���f�L�1.�D���Д��V?��S���`"'�1�������b-s��k*VT�H��D�(fAx�R��!���]�����}߬�i�1Cx�<^ 4N�|9u����?
���T� �D@��ϖL�1�Z��O#�~

����C�2Q�5��w�a�=�}�T�ƃ(o<�8�:�h�^ms�J�������Z�Z��֌q���60mDwޣ��M��?!:�d��1|��r^�f�U��Zѝ��:g8��f�0�S�*�.'�~Y�^��&p�k�w�&{���i�H�y��OPG�������=*���jp�y�(H��M��~h�݈�t��nK^8l�0�<�x�Ezm�p�Q�a���w:��4��e;�vY�(��/�R��8��/��(Q��.�`&�v�|�R����7�a����.]����M�&�9�x%'q�o�S�r#*�{��F�er���D�^�628�,�9�|[�x�rpx*$���.���vB� N^J[�̕3�X�7��N�o�<S���m{W\��9=����V���o�)�#�#]��m
���lP�%��=�_�Þ��(��dHstA�j�<��t�-�^Å�#�|�`Sp1K��K�ϭFSO�MpI��ŧ��E���mئ2̓���t���\�E��ɉ�Q�Xe��oL1��4��A����p�?{��L4�;@�P.s��&��\a:ى��0	E������V�@���
�' '�����ʏ�l}H ,<a�@qҍhZ�u-R,���^���+��T���<F����JwP���-|�c��M����^0�@�/D6��tQ�|������G��e��S�yw��J��0�3����?����˚[Z��0_z��.w�Q�_'�H�DF���+^̚�e�:����2�u�� �v����rZz4&�_@]wd���,�Z������H�	I�5S?8+�*��V��{Jt�0����^�9I]u�K!O�n���ΨD�M0� t�d���5P-��e�*U`4�w���y\'b�Ƶ��72_o ur���vM(A���AwL����@ߏ�����05u�g�ë n�$��Yf�:L\�s�e���Ksv�܎0�ՁL�ufٕ?���26u�Z����v��_ ��-� �N���c��XT�9D�0�Ϙ�5�,�Q8*_\"��Rc���h��tc�&6�Z�cf#�����30֦�*��
���7ٹm������1�L��ώi������f{X�V����3�����e�ǽ���'6�%j,4
gT���t���_^�~^�f��QR���Wu&�'�A-�װ�WQ���bM+<C&#���Q�jQ��m��Ǚi�8rv����n�D�g ��aa����-=�(/I�K�$��;�V�J�3������� � �l�ބ���¯m��HW�8��~xZ�5�
]��d�-w�%A��tɉ#	*�&�l�'�Rt1��^�դG�
C	�+�z�É���l'�ڄ��	j�C����3EaSD�,�Ƅ��6�L�_��j��0����"�$�4�rЅ�]�ߟ����@�/d�70�D�Y�u��xu�$�/N�w��Z�
7��ZX�,ܒ��=3KqT7c������.��,�:l�ϔ�T(�>a�
p��Ϗ���E�D0�M��)"���\R���[H��|z���*tT�Ж/ç���@�B��%?�.�D��dr��BA��&BRZ�|A�\	���=�Zx�C)�����6���yn�N��a9�/v��r����e�� l|��f=��
�v�'��b�զ�J�iL���� ��#�f�2���C���(۝I��������Y��i�nk�-���^�K (vpf,v��gʙ֯�� �������-cP�i�E�ò�ST���Or\:�js�A ���E^��{|v���9Qdv+!���6Ut{y��~ɳޞ~�]�3��!����z���|H���q�^X�p�NI
-��ĸ�R�% �9�ƿ�B-��[/�U���G�m�(rZpY@�C�Z�ǫ)yh ����>�����9``�K1 ��%���7C-��!�`*�f@�*�6���7MqU�f8���<%3��a�-�7��\$���@8f>��@���'�U��8�8@+��@JLǥ8v̙�p:x��+b.�u��<ƭρo����`1�o�+�I��~�]��M1�*#��H������p,c���ZD�����45f�Vt]��TVYsc�� 1��"cי*��C���ˎΚ"�lO��2�6�-R$�EޞS����B�Thɷ��jiΗ䈴��g�F.���`f��'��%��a�{��>bk)׀Ծ�B~�������~m����.)���9ÎuexX1iYɣ�����=��m���8<���4��R�
x	��?gUs=ұ�\y0�1�ұ򹮷��Ty�޻8��]S����~�ԩOwj��&��kz���Zm�s�(��!l�=�./`<��*Sh�%+��
�l,�(pre-#�O����X͠���]X�>��J��P�+�m�p�p#h�EZ���[0g���B��&B�����)D�lɰ�,�<���1�1���Pe�V�3&�:-u��@� �aM�]�^�T����}�D�}�5]]r���Y\��bo�y�|�O�1��.�������Hi��"����y~�-���"Nk��1�o40)�-Hk���0H�`��nǞ��6��!6�z��ޞ"P��O��R ���F�Q�6r�Ez%�!��k!G}f�o�q��&�~~�k!@}xaH�&��h����rɯ����&i��c�UEn&\�N~σ�5h�1
	#M\�����tUC'�n��J��4e���Oj>�9��;����Q����x����9�߭�cQ,c����}z��*��,��0�t��H�~�t� �[�<�ϴpw��ɖ�/���H%�zg���b��,)�.�ى[�%i�6��=�3���q5�*%$�c�n���+��t������Zh�A���<K�(>��;�p�ͩ�ؿ�d��X���.%�v���v�X�;Vcm�]H�J��F��;�+�E�<��evƑ�,��n�� ߢ3G}e�ڥR^��sS\f��)��-#��*۵v���0�غv?����N�D�8��gJ[�6������qDS8�w���$6�,�n�h7�r���]z�hS�\ݯ8A�^�ݒf�96~I�.!`2%��q,z*��e<2�uK���j�m��i��5�9@�P�v�
u�~�d{~�+��=�*����Pz]�G`���#H=Tn(p%�R����^d%��S������m]��L��
�>B8\�0_'�%����(��j�o,e���q,'�~p�^!̷xş��(�`f�bβ:&���pB�	J�d��h��d��:�b-�>jpbXಘ�����.3��Y������%-�A���H�!zFJ?_w��:3����rg|Ua��q�E|� ,�RXj�g�d����M�$����}f������ Mc���h��� �SK��v��\�'��A�T��F�RJ
�F��,(Miݍ{���:���>���ݬJe��7tʠ�["T �@3;n�"Je0���VRop�|/��ӑ���
�ӥ�
�v#MŦ1�)l��PŖ��P��Jo��W�õ��D�SS�{�;I�`�OM!�Q�Y2�ń��?N�|��9�&����z*�d��Q��q0�q�Kg"��M��uOR�i1���/Te��o������ԝ��ͭY���yY�1�2�c������N���劘M��U����y�'H�y�a��qՐM���$-��]��т!����d���^t�u�ٚH��2�0m�dL�d��}��?��h�ᦷ?Rl��I'���nıuB�Y]�Cρ<��Y��#��fi'���"��*"���z(�eF�<�\#�z����.L��r�u��?uC���9Ӗh��.�s1m���6T_����r;l>������ ��gw{E
���Gn�����RJ��bDC�FbU�L9�J�e�w~�"��qԀt/��r�Ec���NB�xw���a�<sa��BL<Ow�#C�yd9ӭn�.|D{4����H�|�uX7$�v'�AL&@��D���@�"olx�,���d��HJ���Ō��7�*אZI &?/�I�����[J..��o�S��)]o����$w�G��+�r,�>v��
��LF�]!���:o��� �V �FP.�����B`釡�^C z3h��I	^T�#&�Q�p�-l��_�`xD5���w�v��U�ZǠ�,a}�&�	.���F~ڎrGn�7�)a;�S��>�(�:��E"q�\��"�w5Ӻ;���R��澻)_rH��^�8t��?�Y񡀋N�,�d�9(t=ä�_0�i���ߐ�t_�EZ �9��� ��^�9� {=���r&]jM��83= "Qp����=֣�¸bf{V��ı��s��[��~��49m^BO֑.��&�m���Rb���g��-D��&(,�.md ����p,O䏋�å�[#��h� .�&��/8�LxT?�8��|j�y�ub0{�Mo8����]m����D Y<��;dbc>��j|!D��>��qI�P6 �{'~���S���F�k�h~�&�s-ؒyE<*H�X�g*3�`p�YY��m�0m�����^�џ�fA5p6dH�19�ݏ(َ3M�%ހ�rW��e���皼Xr
�;����gW�Q����@X�c����:�
��t"����o���)"�;0~o�H��E����UЭ}k�s_�n��h���HAM
�$��5�ѡa�qԫ^u,�>�DG��qO�$��;�b˻M�˧��ŋ�=p�z��b`�b��&�/2w�]@XJ��R��7�
�Z�4��#�a�5P|�S2�god�l�UCS�@@�ҫkg�W/(�͋���M�� �^��O���u�fI�~�X`��1��\n��	-�)G��$��O����`*gHT3�f|�B���*Du��Q�cJW5,�����9M{��ņԺ��_ŗ
h�oG����@~j�����P�v�*$�a7�#��Ld�Y���+��5[�'�+��KD1%+�첻���UgJ�6���;x��Ư� �	[����:�֊3:�	� �p�@Ks���5�hV�L�k�/n~Ǫt�ս̣���,hy�r@V��^��n .D}`�丶���hc�������k�A_�b���� ��N�r�{����?	rҥ�XH�<	S�UHE����J_��G��d����ɲE��%IS�ϩ@a�=8�T���(h���+�?=��rHٖ@5dd�d;������>����@�jG�5�J�:��v%��|��:2�5W�~&UXb��;Ѭ��傣�+�	ٵszD@�ћ�Ш�Q�K�ۅ�>��2�D�}/�\
���Ҁ�W}l�����#�^�nE_x�bf�X��(��47ԫbɔcV�R���-Xi׊���S����:C�O;�
�M�QQ@��(>3z�f{8���9�8�����l�QؿJ�D���]�G�M6b4U�d�I��QMW4@�@����銂8� ������i�n�・��� F�P��.	ҽ"���p'I�jw`�HQ|S�Y����{��H�jj�}�Ҿ�gKO�� Y�>U�A5�D+z�y���|�z�ej���v�}rw���k�t*�(Y0�U�����`��&/k]!���b-;���W��ʌ8F1��a����ߝ���J;���_\��� <�\hu������V]0-i};, W�l��l�i>Ǖ^i�kiK���E���f��Û��U�`�M��s��F�?��Q#�܎�qW���Q��I�Q1��\�?+h�Ubx(Ds�f�f:��\�P�-$Ŋ/���
��#hYw��bY��4>:����[��O+���F��"�B�L��#?jx��n���.��ݯ�^��F��#QcI���w��w���6_v���yqG�&�US}���ѱ��8��c���-A.��dWޔ�[�x@B��A*n'�-{c`+_���0�\�MOS)�^H�
�h��;cK��j����w�ϲp+CsO)���R���ӊ�D��mѭ��-9����h�b�5��{_�yW��=H��q�(�C,�0��ۀ�� &%&���w�l��%x$�vќ�Z�����\�Y��Pl��I'�hE�!{k�� 4-���v����/�uu�R�#�=R����=<U�$GQ�<�ɬ��Q7�����K�3��F�%N�j��c��;�םR�ὖ�ʦ[�YL�����My6�ť��B^|�)�zx��E*d���ݨZ�X_��y&�����Wź�
���J�+�l����Q3��0Q��r�)*U�m�4�z2EH�.�o�����_�G�4 ]K/�sDpCQn+`�|�����M*��\q��G�iN�w�\i6�ֶ��}/��q���>������5�u�W�N6�����+�PdvΆȬ�^�	<(�ᤣk��Ji!6وXZL��|�16؁CP����d"6���39D��s&��nƚXh�2��o���WQ=��1�jT��dJ������7z9N�e���3�=�Y!#��]?��G�lX�ӏ+|�Ĕ�R?w�#��~�P��͐���g���r�Z2�}��L�1�5�t7�>���}��`w��({{����N���W���ԙ5\w��4�J�E4_0�����_�ˎfI����zNp����\$m8k��Z�H�_�R��Β鳞�x"t������n�1ae�Y�_��8������e���XԚ��{��w�6/+���/L�{�J��k0�
!����:e+�*�=.����M�:j�5��W䦦_o+��XF��kS5�ӛ��*�i�7I$WY��C��Y���˞l���I6�~�e�2>Prɜ�gU�~)�:er� � �d���)�iUBqEc����5� 嬤�����6ġ{���Vj�k;�L��I�2��K�b����*�\�f߳�)We��w�I��#�y�I�Ȗ��S�^���
��%�~tmrИF91���m;�#�GڒZ|G)�F^�W�����	
�|�?����P[���"�H�Fܝ��\�#vVAs���R�1N�=è��5�~������Ũ㽯h�s0������K�T���;���Om���u8,*�zH�Zt�F�3�;h���X=Y��˒�zٻ�%��Z$H[�ǊL�u�B��ݶ�A���U�M��<2�#$��)'���y��3	�u�B7�NT}T�iZ��ovא2/�oː��x�mZ��� Ѩ�FfV�fE��@�<�Ed�:z���������,f4dRK�';I��Rg$��6]����ȫ˟(�	[��r({�� ���%"��ªW�ȶ,�e�r�T���� C����Hɳ�#�u|��L�t������Dn�נ�a��o�a@�i�n�0������rL�_3A4<�����@k�����
���H����˿��-��z���yWm'-��h��G9�7U?����!�@FJ2�3�f��g��s��V!���x84��BǸ	/)�b�X�����H*��\���	�<�%�Iҫ�3�GH������j�KsS�)ǋcz^u'9ٲN&q�a"w�r'��[I�c�5�u?2n�{��DQM�⊵kr��@m���I�����=���VV&�hI��3eJ��� ��V�Gh���3MĎ���� #�9�'��Q�jk��$&h�T#���տ��=c���&'N����9x�kg<���C�4�hs��b����B�Cv��k2߀Rq-s�����Hu1�.ȣe'Ɩa�bRh�/�#����<�J�	�A�f� �v23�e�l,��ύ�.���Hb��b�؅�*����1#/o��3/�WQUi�A*_q��m��.+:|[�,QZnޢc�1��e��V;�+�P<�@�˪P9��n�����Y���*�����~C��ݺ�v5��{6JE}�G��X��_i4��f��0G�N�T��?�Z[r�H�2�^��3�;��t�B�4)��"1�W���v�1��Oʭ��o�&zG�d��V\����'ʿzMЉ-���5�٬�i��>�S�>�����6�/ ����qlvV�eG��<���Z�*�6�\����j�k���&�@``��ڤ���&R?Z��MUZm`Gn��q�ˍ_5�n�0]�$&$eZ9I-����������Yoq`"�)���F�vw��'��4'bc������?��aTh�C$��@� 6D�g�JP�
�j�����?�	�NNU ���Tr�,�?���B{����}+����/C[�
�-����D�uz��v����=�B�|/՚6o����мE�-
������n9-N9���3�����у�A�D�C��%�j���lcvx4�_��S���b�3m�"K[8�.�����8�g�;%�$Q0�ʾ�YΨ�Ha�N��z��|1Шb�ԭib�s�曬�E�C1���I¾}���q�% �R�:R8�T+ŚT�-V���A�$���Kr�Q���K��N�rb}��0HI0�	͹�Z,�������{��Ư7q��?D�O�����X13]��5;-G�{���h|��ԣ��������os�b��Tl�u͘��!/Z55�IJ\<pg�yd	�;6�h�A���gnڽi�.����$
m�s��*�Xp��ډ��:c�EWשPO� $�'"Tkb�E���'0Ҟ.*q�IR�׷��r�!�(���	+-".2`��R�D���&�B�<AA���C������~���J��9-�"m��b�2�CΟ}�%br�'a�����!��gU�؆�� �׻�1b�h����8����G�RwwEH�����P:�r��0����ܲ�@9�n��*Tb�蓜W���v���ÿ��<�MJ]�aBX��A��Z������r���)s����b�GX8]=�y��1���gӮb��"x�
�0�*r�ј�\�Yf4�l�R�I��*�q�(�~��u�N~�KXl#{��Z�\�Ǘ�>�>��#ԗ{݃WExlx�s���M鲄�?�K|��ƀ��Ȃ'-ZS�ր,gTַ�a#x	3'2�z��<��Ą���r ��t��W�t�9�
�����m�@��C�I�E� �W�SA>��_��V���phx���?���w�1�ER�9�HiD��ieu6�#�˝�[X�s$>�-z� 8ֳS���7h�jJ,P�k
��X*G-�?4
��p�(����5�<o�9Ow|�B=��Bf��0xw��R}�烲�&F军��10����jM������6�l�(�'2�۝��y��e�)PW��}��Ŋ����bʥ0��M��4O
ܩ1n���[��(�^Ī��&ߵ��4��꿅��=�����%��J�����6��u�?�eK���7��M}cVR��j=R�ړ��^�E�d?O�]V�o�}�b�"��b��¢���Uz��I�-yQ�&�:���ͅ��&7�m?�z�C�t�#�#�U�i:F��r��bՁ����RYA�<0g�<ѵ
j+j�bD.�^��W5�g�t~��sn�!3�5L�W�)�F3�J�f�X��~Q�\��V[J��)�.yy��a��B[����{�J��0t����Z��x
�����;Jb��	/B�2$
pa�dX��H�����xp�&�j �m�9pPRf�,�P�q3�L?]�a4���!�fR&�0�C�y�^tj�Ż�;�prS�F�Iq$&;S���Į�����������H]C�i'ud����6��X�u�*+��		�Q*��9���#���ý)��*��\dI��#3�e�ݡ$	H�����6,� ��@^>{M>ުZ�/�����2
���.$�"�:���!�´������k���60!�=������B����(��4���21v�]G���5^E�p�s[gsɋ�J:i����M^��[8�kVL�s���W�ŧ~�;�p�R'����F	B
�f]�Y<?�3�)y����m�;���o�d���� �@lN~���Z���p����u��^{�9H����p��}��ƅZ�R5�~+KŬ��=?y�;��-�u%	0��=�.d�1�H>��0��SߧqO?W��|��>���k[�3t �g�5\ ��bh��q�y��Y��3��L~6�`v����{�;�_.c����1Lg��g��0L���L����h.����nC���ժ9��h`ɑ&�_.+���V�}�;��O|pɼ�p}Y�8b�an�+5ii�4�8�gӄ�w���ٷ��n0.?#�֔�J��곿��D}���W��t>k�u��
�$
�Ez���L���i�s Z�%����������7���9�"^L�s1�d1m>�WF��g���OhG! ���Ų�P3�e{�@�3�P���DTJe���JPނ\k��Ҫq����3��Ew��T[Y!߳����1TF ��l�5�4QghӜz��88]I�r��	�}ī7�@~����͸����C�����V��^@��p>q�]^�luI��Gp=R��%8���EE�g������39B�����en햃3ioOz��FM����t��uN�[J���vrD��1BR�z=s_�BnvV�7C�Z�"�Z�X���h�p��ܩ�L<��X�:v��!fټg�����	o�͗ <�c,���Ό�����9@��C5J�	��NJ�Ԇ��EB���"���VF����o�4�M���q�H)L	,/���u'*g�fΜ�gQS�Nz�|'?�w⼆���:'��J�ZOu��I�^+��	��PV�����a��&�ŀɸ>lJ~H��-�);zI˽[�S.�i~����=<���n�_8�@��"�(�-:K�D>Wd���f�+�4�o]�m�����[��Ct�0�z�ٕosz�������L��>����B�:�Oq\�R1��▣ԃ�	*+vF��P�Ҋ :����Q�۷_%��ܡV�7B����8��Aײ�ơ��xr��.�
R*�W��cd�zB���VC�&Q�9�fc/����rg_嬨S�[������k���PjG&�|0c5Q��c�_ Z��jlϪ~&nj}�&�RI�S��Ea،p�6�2�u���=���ڤ̂�}��l��^X`=g�nG��ڪyR�na�,k�Z����xb��(�.����	C���-��ΑU	� ��s�e��|?������3�&M�s���fJZ�8����i��;�K�:��2+�K��k�F��D&�-��{w���F�+5�����kZc�Z0N�:���aP+���졊��f�� 2)��
�;ܸ��L9˓���Ց���B���i��8��/r3��9_�pFY�P��SPk�I���w9i}������r[���%�f�U��6,�sLI��
#�~���=Qe�g�XE��a��@�(�V��� D�,N��J3D/m�;���A��E`B��Щ$ ܠt�^�8Yk�6��(�c�����*�8̆ɅH�86�;�ࣖI�!��FŽ�t��}��l<8��;�D4�)A����W��:�?3��9������CU&�z�iIJ�6�j�X����>�:�:ҳ$��D�t��#�ܫG[T�q/Y�s�f�H���4����<��`�r����V~K��I$�ٳ�&����e�$�͖QJ�u`�5\T8&X�v�� ����p�;���V�i������V�b
�݋U@��?�������3lk��e�](#�`(p|��x��^�P
��L<0,���Q*S�]i� �47X��֗ehϕ/5'�b����?��7��b/8�L3�LYYd�m��F���	�:\[�8t�~6��kF��Lz�u�V�,���F����ɇ�2i�?i��?ެ�떭�خ��=�K�g�t��DN|:'�qb�� 懛CL�����ѿU,���,,��y�!��]� �{]����_f�|{J6�s�LT�u%����I!�u���V��9/�����QjF5�3b��L�!��̽�{�*�
L�R;�������J��6�(�R�^��8�OM�e��a�8
8������u�G�E �b/y�'qN#m���s���ǟ+�)�K�'��J��+�)�����NG�����:݂F�3]�Q�_eL�]�ʥZ>�cV`1����.�Ί��{c[�tj�P{
sc�AK����i�l��~E���t�E�]z��l�d5���2��@2r��1�L������4b�ʑ.���t�Omr*���{y��Ц�(�ӗ?�k��Nh�ʌε���M5۪oŗqB�&،]a�yf�M
_��7�t���P�^5~P��+vZ�?����g��SiuQ@�]]s���@V7-6��t��波TCG�4�{�o� ��[Z�Lğ��S"�!��o;W_��\��s�In��͚�W�0�0f���q%�L�����"{z�D���d�QR�%B_+ #�zl���t���Fۄ���}-؆<�i_]7�KJ�_�,��U����IV��_���3 EQ�u�����Q�
}lM�6M�IF�0qt��d_l��!l��x�0��]$�.�"����LO�5���*���;p��h�����,V5cR{�l���F��
L��J+��L����ǌOWI��jJ���*�,K�B�ca���~�M�.���G���)���5��iqI~��C�xe�F�3���>J?L(4���	�VV��{W��xk5L#G@YDA/��cʱ �~�McX�����Ҏ��s�G��N2Z�Φ(zy_/p	�(3�g�_��Lh+&��K����no�k{Z�2��u��}��
zӼ���^G�w١ ��.��b	#���ٴ5z�Ih>���,�>'�]J��F�Ɵ��^���'c
��M�'��ݒ�(P$f#�t���Mj�Z�U�7!ܴ���'${.D�s�4-�2��l�Mk�� ��}��7��;L�i��ը���%����D�i�w��w��"���r$�T�`�vХ�k,p��7��_#q�ŷ�C���H��yXzG��D/<�^<�����S@�b�Tq��T"���j��R���b�ď:�J�=���Y�?��U�ל��;�tQİ$.+f���&�V�Si���A�a�xsԖ͇~M7�?g��I�q*������w^�F7�w�z~���l�7G�מ�Ŧ�*$;%G��/�d��ͻ��f;��7��ÏA�\���.�*�K�Y.����v�S��b��A����C�2�gs���ϥ0��������H#�>�I�k�?,��n'\�>e�ի���B�ǉ��џq���<S/�u��t�q2����́LӦ$(T�o�s�H#�%׮fY��eYJF����t�e����d�7qЕK��3�s����,�ƶ���ȶ��Z�o�!Ċ�6���)��~��\���8ъ�,מd]�Z{mp�K״�g�q&I	O�pk8g�(	z�v�(yh�G��g�Q]�N�N��WE�0Z4�U��&ǒF�F������41���Z �5j5~g����"?��m/[�FW�CoVp����h��l*.t�A�E���C�J��s��_Ē1]�5�N�i�Ȉ����r�n+�Ѥ��<ōh(r�^w�U�.v�s���Q�o�AA�ˤ�	�$�;�J�G� .��O�,�߭:Ӫ
 I�����p3���"�x,廊�Fɥ6��=0#k�&�k;�Xn��i��u��pw g; }�mp�agb�s�y�+Ϝ�t$��'��v�m�"%k�Na�.�qُC�<�BS&�C�.3�"Y*?���f�/Qy2�[b#)����*7�gOB�_���J	�4�4#��g�M����ωQp��Mt��rI�LڞѸʒ/�P?��2�
���<���#� j�C�0�^g�IY峎����ߚ$�c;��&��$ߖ
�bI�nq���ҝA� *iFғC/T.:�� )�-��C�T�x$���#�pr���7��+CG#nm��w�-dv�00L���qn!v�Z�W���:4��c��	���g�θ=�豽��Unnۘ�:~�3?���	,�r�*��.̀g�Sp�m��1�˼�5��FSy��e�����{���&���=E���ڕ{�p��W`%�0�r�D��ӗxFKϟ5̮���ӵ_�(�k	��@��$o�(����t�DS��X�^S- ��i�e+ׂjk7����H|�����M��Vw!����e��C?�V�E��&��j������k²:Io������|�������1k�\�Y�S����?�?�?����\7� ��7��5�_����x���Dꃄ]M����hq�{���O���x88�t�bY#m9�������`�ip��k�LىQ^�Dڃ#/|㒓L%bAy7^�,���^
��v^��*���j�D�KDA�(��DkW�ި)V7���o�G�[�Cpv�C玵��7Q��7ۭ�v�5��M�r��>.��8
�cx��<Z�y}J�S���e1�U�*���f�T_��&���0������"V�z����1��A���Y����Х��	\�m=Y1��u�.��|��\j�#\�]{ �z/�73��-( Ti��6Q������ʞ8��^��5o�
?�j��n6�o�<.>$�R���{=�)O��{Q<���}��6��SA��l�����몒��޲H�dIϩ�i�;�ײk��[��tW@X%�bŢ�Q�&v�X�dd��g^�[�FO���A#��1m��}p���`�`��R7������J��W���1��חv�TE y=�fvNq�|�e��Lz�����t�3�+�@ǯ�F�T���pk���~C�5��{va�+1M�N+L�]=}��ݝ+d��)����DQ疪��������mx!��hS�˕�#L�tTb��!:gPw�&��]-��-�`뢲vc#�R�m5s��9�9W=�����OXu/���o���(P���x�\�i�ڃ��g���?�r �muw��/�����ݬ�H+���-�� �E�8�[@0$�31F�Y1���w��`�h�KM>���3�^�Z��>�
��YX�ʏE�k��U)�b[�(a�B-�ii"���3���
3R�v����:�i��ኃiv�Vp= f��uׅb�� ���	#��)����C�y��	d�|4w�B�bt�p�ԯs��X�/ݹ;�)�g��Σ��<� P~��9��Z�/�ew�Up/�2�
�^���R���� k����I���-4y B^�8�߄�+�F�t�l,_p�^5*�f����w����;��\a��1��E�"��_Y?X�Fm�l�i�c�8<�j��E�V�(3\i�c�O�R�l�@�����Ht�n1$I�1��� ���������J����E��:�_o�*����/w���D6��|4��\��1�P�7�"����"�@u��ܻ,�蘿7�B.Y�sp���N	���%/�~�S+��q|���B\'Mt����/�|T�<ơ���03!b�pfX]+�1����zL���PCA���X�2�	�Ƕ7���]]�&1����4��i��|&�ZǇ ��\�14�ʆ0��$�c��QM�M�Ę���Uf��ѐ��[��a�D��߶ړ�<�������ΐ�(b1��+��0����M���_�$7�����X�Ôֹ�ό'$�� @
n���vp�K�u%�s�2��#�.����lv�4�B(Dh�1JL/"M?�jׄ*ҕs�V�����wW(+c�[�icMWQ��ꃧ���O=N@�Z�)a'rY�F-ŞN���r"=�fŕ_�m)�+�m�2R�bθ��N���ަ
q�W��s�Əis�i
�+Ÿn���Hq����7g�R�+� ALa�X�����CG�j�F	'����GGdF�8ٞ�l0����&��0,�`�[x�� }�U�_��B�M��CG�t���2�� 
��G�p1�����'�`���o�ĕ.Z���p1�����9f�\�~�����`F��|���pUrI����%)��$1��Oդ3d�.��s��c�~�YI�sR��ۈ׃�R	��������$��m�Km�5��p'��uW#���H��_R��%����w!�s�o����M"������|A^�6���>�U���ZW>�����>m7wvm���l �	
Rh�u.�(�ľ�Y@�@Uh��"�tql��!{�R���&��-N�Ƥ�%?�]���i$�j6R��ˤ��CQ����]�Wr�`)E�%8y{��W��l�i �c�d��Q�`����0'�;�me y~�fe����*�˔>ؠh���]�Gwȟ�5�8ƨ#�Ƕ|�~,��d	�K�a��\Q˘�iKu�tG������]Ku�́�_X`'����
ye����ܬE]����1la���:9d�k�Fp�C��I����'���IͿ�u�E�i�ؕ�8�x��lc^����_,���t��,�bh����;m�Gyju}����*�סf�3���+�R%�y���/�q;��2
C�����;���=|X�|������q�{\/yo������.�kn��e6��B�"����'��5d{Բ��gìC�B4uK����&���t_ ���Uqs�_��!W����X�?�X 6��Ǒ�m��+�նm���!&���v=���a�4v9�B^��W���p�ţOt%$g[ey��҈���*�'
����� F�O4� �bn��V��/7�G����������;�u��,j�Ij���_߬Ҏ��1�h=uSg�%=q�j��9#X)���nb������gH�!7�QǍ�/���R5w;�$���>svʡ��yPx;�pĕZ�7e?�X�[�$�+J�����Z���k;�c�ҎO<��:���G�;�-�U�s�K5�Қ�'�O�aB�^�?g!��gc+7��!���p:ͷ�d@Q�JRq��u���;$M@Rz�~2>Or��`1�( ٪�Q���Z�uN�D�>y����D�,�
�"�~@�]VY�a>H�i�r	" �� �9��`�<dJ�>��b���d�tr]q�7pO�?A�Ƹ��[:0��*+2�
��r1�<4���Gb�g�QF����j���T/b�D�yN␛�'?�b�������|�`WM��CE}����bɮħe�M��}IQ����Q̾(�~���i�>Ջ>�tIC����[&zW�����oq�Fc�} =X3���"��P ���
U�t5 �BL�C$����Fyឺ�wv�t^l�ݧ�7�L1��V[����dc�����	��P��y?�d'j'X��� !s�:�BڍX�|�!�0Xh�`��,S<�.����H:R,1����oV�LI�z5����i^�9�׳��W��\�}g=}d�[	r�z,v�q�rƸ��:Z�
�N��,<���E7h=J�ɚ�H��s/��٘al�4��~	FN�X��q?�DL���M���@��&�)N���I�ë-�����-D���´�'�T�|�_�/,D�gO���p4KUB���]�do��_��:��O�diL��j��v|#Wj:*���.@ߕ�M�o-5����Q���3xa�ȭ1f�|�E��u�a�ϓ�.!�+Hψ���}ŭn4��O%w�f=~p��P�4#�f�N4n�⍢F�H��Eo̻����
?X�L��B&~2�'�Lj���U`a��I������)1p�*���(�Tw�/��\{ 0Ú��A۞�=P��Zg�l~F�6�|~o4m���ػuri�0����"U�'��XRT��BDh]�mH��$�����E�[kȒk`瞈jG=�8�(�o�Wy�$g�*����j���	Ҍ��M*`.آ��*�k�<#�t��&�7$��	K��l��X��u�*v��{�_&۝�_I�h��hi/����(�t� BƞvZb��mڸ;Wb�v�߸����x���0p����S�Q���-��n�ej����9�us�E�˸
���F� �����l��gb�؇e��Vw���"�dj�.��4�@�ȟ��=q:,�.��|�=@I�Z��ı�%AU��#Zq*C��x��I���܇K�L����
�\�m���A��x�%D����n�K�Nt�!��/䎂�:�q�}~�,�;��N탾Р�09�Y1���hRk�{��>�r��0e���iA-�u��1�YAzemw${���ɂ7.��iK�Vm�3��w�O{������	�����cJ�4�r��)�ZlA�[܏��s&;�����h럋4-�(`��<p��((0FI#m����5�HS������q#5��9B�u��3o#�<�}�"��ǉr�h���8Ϝk�I1�1
�뱪se�l���ɪ��Fw��8��'���drb }�rv6i�����:Gx)TSF�hq���|z*|��x?�c����,�,�c�:�yF�h��(!���i���a"鐮���}>�Ʀ��%c��ueQ�-�����sr�l�b^솛�4#�)���^�w���^�{�HQ�{W6��_ʑB����� .� �c�;�es3S�406R�_�ڠ`�b���P*���Ys]�[V�,u����gT˒�ǩ���	����0t=�`�0/%�^B�4���F��{&�"���Ah|��8X�ߥ�:���C<*�ѭ�\�_s�!	����U��[�g�4�R!>,T*��QN�pw�٢��-dB!��:eG�(P�-�� ��+c�Ĵ{����R.�mr��1;�P��}rr:�r'�rL��zA]I;�Pk�Ҿ��ʗ��T�P�sj�>�>�kv�)͑�D��}YD^�/���t�:�ܹ�놝@�̓�87亴���`��=,P�w���W��oY�W��t~T,^��˔��W����<�Y�4�64���) c�x�S�4�!�?����S���/��'��I��Ye�5����;O@�=ΊMH'���y@�8&E:P7$q%��@�I9-�c�����Vdg ���rhB����VCZ�1�B���0��fb��l��u��@���-Ki1]���H�@����Vh)�h1.�N������.sD�=�"8N��T}�[�3k/�h3K����\��
�;5��Il�O�uJj��&nDcձdZ�?�?��E�_<���}���LUʤ���y��$n��!�
1}�lUa���:�Bچ��*�CZ1�/���(�P�/��#+[G��@�$B��rQ����d�,m>5��Y;:p���K�����N�MH��nF��-�_�Nth��Ӯ�H۽_'���N�c��
��*P��>�c�wk0���K�.���"���6>$9��{ȘJ���izH�*	o�1r�2oG~"X�djO� ����P��Z���3��c���M�$e����8���{��l-I50פnx�!Q��x028��E�S>%n�k���V�dN=zK��mD�i���:�9��	u�y�QrG����:��m|�9h'7���]?)�w�5�q1R��*+�rN8��ɲ4SE%sy�v�O[�;�@�;~��.�:=ס�_i�ۓ�4}��'��x�Q��9%.fsw;����6g8�Ԉ�.!�n�>�s	\�X����y��̺C"O�n�]߸���n@�9��i�ʇ
�S���z�G��\��UQ�E�X� 2�k	��DHA�Ev�*B�|�1izE�C0����
-cn϶����Gr���U���	 US�i�Ύ� �gF��`�ZRé3_����-��axQa�r����>e��s�"���	��*���[T���F�mh���n�>�՚�bq�9�?0��ϭ�n��C6*3,�<��9?��f��/��._/,�ɞ(\;CF��phx��C�JE$�<��MW��[1�iF�Gw�"���(~�@ћ[Ig�>��<�P �'YA��k\���꣖��*Aɪ��Ηn����0����]6�B��$Ւ���/Z9�|)dJ����+R�(D��0G?�4 D��.g�C�$�-�G�.��hO��ۧ�_ڣL���|f{nj�:���q���jOn?�����m�Q6�*ܶ�OU�=���>�[->����F�n���B�>�'��X6�&�e�k:Rv�M����=@�^%.�}�a�;@�����F7��꠺pG�� �����Y6���	����%Q�� �C|���<㬄1LYJ#��^Rk�U൦���]l�;�#!�g`Fk��f��K-Ĥ}W�oepGj�r,b��:��{�f�8���,�x�k�7E](N�u��R|��?J~BrI j��1/Oø��Q�����<ӵ���a�:i�[��PکW��3\�{dl��=�����uVC�yZl?��Z`���M�{إ�̾����t�I�{%�J��c�uL�\yf}�;��r�m�����E���������L�t���v�����Y����s���{�Y�w�)���?��G�}䳭���J��Ǘ�qF,�M�η�g��	(�n�J�8�2�0�D�'i���ܝ^H@�߅Il�L��B��z��j�����`��6�C(��]�Pa^!�-�B�����SY7�Wlx�ֲ��xN�#B�T���%vրJA9��������$m�a3�V���g��P�&�۱�w�Ɣ����>y�	��a�4ZX4l5Ӂ�T��Y�~����X������?g��&	X��N��@x�P+��/r۞��%��z�ͅ�"�ԇc}v��|z;٦�6)Cu7Gv{i��c�֌7̂'�4�����U�[��i6Y!w=ۛŃ�xQ���� ��ek.2Ją����w=0r�d��x�`SҜ���~�bޟlH������^��
�~����A.���T��S������q����i�,�VfK/�PM�7�ˀc�Ꝓx�	��VVI����j@�����u89�_�K�L<�|K3���V���Uo�#�a��=Ȝ�3j��R\EĻ��5����Ҳ��(րf⻾�^H�f��N��'[9n�}d�np�Ĥ(yb���D�[��ʬ�h�ݬ��fH�����z�%ʹ��%�!/���TC�N�Q��Dل+��.�!����D������Ȓ�UX�����#�	�@�2&�x��R�!����}%g��&�6B�Q�5ً�����Hct3��u����i bjϛ���&�K�k������3��M꽨c�I��j����a 3$sZE4��O����%�@Y��y�WL2�6���;�i�UxfS���s�gj�Ź�8Fa�C��5�3�a���q͜��٫��c<��Y����F>w兺"��xS}&<Z�1�$�k���E�L)k7:�E����Q�avGsPFN�օ<P��l��>�.�wv%��;꒜Sm��ƈ׈$�2Z#ܕ/���5g�X�v-��xݢ�sq��������w�r��E��p쟪��[�IpQ�,����)i�+s;[�Y�N�p��!4�"�! mQ�YS��y �U�4�
�[�Y%T$�r��]��T駘�:����^nh[����~�`Y�'`��P��k1/e�l~-:16#�� v�B��]3Q�(-�kƅ��SP�Y�rOA��w_�&�2h��IjgS�n�q��(T�QD}���&�?�g��3HK��`뢨�e�̄Utr�7Q#Z��z�����M>����F�h�'�<��ͅ
n^ 93'b�D�Y��O��LnnYY�:a��q�z��@���Ͷx��Rz��˓+�8,^� AӠ�~̑N���� ɻ�BU�T�@^��)��k�<�@2U=#�.��DEL���n�e6W�P�,hL�,��P"x� z��[��:W�ዦ��*i���G	�;�y�еda��g�95bm��;;e���"���c*��� }t��8��8Mҟf~�W_Bd+�]͗c�e�7���MXb��Nc��PN~C;�֠�s��ۯ?�\Tb��-/b%�ɋ�%"�!���R�dD.;�6)�:p��������Mp�~��H��Ѹ�^���!�t��'�~�^D�x��ÿ�`�š.���(S��'�/��ڔ����^�����m󼢫��Ӳ_\��;_F��tC��Ro����;?�ȚUjˤ�<'�l�6���1Y�}jtL�Sh{�bN�d�k�h��OB�zAF8��V�qp.v=�AkUM�E�W������[OG���￝؅�Oq 1�A}X�㬀7	���H��qj(T�۞iK�����&�zz߈�6 �HB�,�6̡��r�۝���]a��H$!ZiI����d�z�S�M?F�Jo�ͫ�@���"��\�ǁ�ő[�?��e�$)ɉ�k�A�k0g�E������v��H��Vq=�ez�8�R� �\x�[��{hh�%�u	����Ҫ�x膬�W��{X���J7 B/aΨ5�֑�S5BQs+���PK�2o�(�$�۠pn��B�bS��t!��2���;�� ��$=R���6 ��H���q�36�7�AJ�=Da����o�F�O#�����=>Ҟ�?!�g�����c��@�"\�|�l�Vʽ ]AsÅ���,Ru��o.��=�8�6�������t���*�Q.�Dt��E"���',>�E���nR�|<�{y��
�/���ߙ,�ps7bvN�yR�a$��.Z��Qp[�(D	�����q�jB���D��*"'���w���4l��)����dCS�����	M���گU{j����Tc� t��ص�c)t���0׳h��O���jMPL����ok��]zj̚_�6��iF���Q�3z�e���t�਺� ����R�L�܎�O�^�9��/�Sa�&AE�~ �o���� �^�Me���^�7�\d���(`��S�mX��҉�!Y�`�%~ܳo�t!6L=h��;%]sv%�_�>��JՓlxC� �*r�:���nY.U�D���e��R҆��l�p�/-�� 2��>�8�9EK��)>S���jP^Жג�v�f��V���d�o[�]�v2�J?�b�y�&�/��	�u�s~8�i�z�.���e��[�u�b��>On��5X)�{�'��"�9���79K�V1ݭ��7������X�ݭ�H����
M�t��h�c�O�MEWѼy�<�x֌��Iј�I<��֑.h�@���=H�K�N�1k����JVZ˒���<���Dtm���e�ys��]�"U�������leѝrh;w�P��iDR��:�CS�3�#!KX�Vۊ����S�gІ�gO@yى�de�wzӑaYF���汭��Oqrc�Z W�Bξ]����VcC-�j�!A��Z�յ7�U���z���Wu����5o*�Ħ��Ju��M�t��/��0B���:ΙY���Ӟ�-�f�P�܌c�f�yÙ���4�2O3���w���h�p���|r��W���i��>/8��Q���3�o~�	`��Q���WzG��SW �Y���t�]١]�hgƄ�P��3׈����3M�_i����P���cZ��\R"k+{S��d���L�w�P�b߱�Z$�宄�	����k�dn��C��tE��UJ�2�Qm�Av�N45���doX��9!<D�Z���rQ@n��5,�n~��P`����D]j̛~���x�i�{q�)��Z���$S��
��������v���M_,uu�cΫ{�����/�d��0x��r��A}>_�s�ԩ�P%�=�ژ˘sPK�X~�½C��Y���Lm�M�!#�6i@� >�6�;Ҵ�g�� �9�m=��A	灯d��-���҉�2��N�\8�Y�͟��O�R Gw�g$������?p�3�����뿇C���ͣ@n.I�Ԕ��p+[�isS�Rd���X��s�������H_�MF@z�1B���a�*�uV1�:��^��3a��;���yS!z��6)x�ė���(^Q�F�8�݀�Ac��S�ts�t1����ML-?$�b��o\��/����m�U�d�QG5�hm��-b?��Q��&�#����Co��IgC�6E�0[�������V���O�������Gr�п�z-9��m�i[���т�* 9�^a�ˎ�U��B��S��ɿ|�"���	��ɳ�_a�I���b�a�F?�O `����G3��=6coyN;퍭g�䜧����k#lGHA@�f৑)�x��jL��#�b�掛r�:�x�~9H����;���a�K���8���܎n������ȫ���'�1�j~��?7���KP�mЀP���EUG����G�}1��MbƺA�N�bՕzw+ܑ����84O}6f;t�b��������'CD.�d���~���H&�H�T�\�f��u�:I��#��;�u�!��F'3���q�P*��2��.��R+A-a�+�p糿7�H�����D�}+"�����xߖ�h���VX�@��k&��5�����ª^���
��W�bG�t��f]��.K��K�� �r4�>Ɍl���F>�z��,�����]���R���\koL��پ��'�g����l$h��"x���&�h�z+6�?U���	� oJFF�����-�OG���?����#7�@�[n��v���c��>��:��V�����I�L�sa��>YP�������<�m��+�t��w�p�Rl{b�2�H��Z�	���F���ߢi�!o;��v�����Bzb��tF���&�z88c7 �W%�B*6��\�X�a�ǛҾ�%>U�o3p�a�xwmI ���o���*j��e��(4��=~�P��s���9��<����= �����B��U�!����-�Y�թ3\�8�2[�Q$��H���߂�2lϫw������,��3e�9��Z�l�ʧv�2�@��Ɓ��C�k\��I���-��y�&�M�C�э�+�^.,�Ų�	WD6N3��v��$�R{{N���z?B��2ሯ�F��M�>'h��D-���7Y��"z#��}'k�`�4b��/�+lir`�R��swO�-��}��$��{�tʤj�'�33�Qg��4�&�����h^�a�k9����DJ�e���L��!�MMpL���-Z��?Ԛ|�MOxO�ӄb~W��~�B���B���V� H�Oi��a��О�Z1k��q��YV	g��.�ͥ�wk�=!�f����ʄ��b�8�\�&�3�X����5���������ɺ���)t�4���.�op�-���pd(]����Q�9f�x�vf-͜�>fIx��R?�2{)�/A$�kS��!��cz�ZD�7�o��]�,�~�VN{�gFSʝ��N5}�orF��`<�b=J�jA�'��6�Rcw]��E�B@�j��+��s��{��/���$D��/�׍rt�T��	6k�0���@�[00s"����7�*�'�氳>�IujH�%>Nò�S�|�@Sh �o�G=y���*���Q���ߵTF˗�-��y��t�f�����@>�luw�e�B����lh�$L9ؼ��!f���(q�C	%T�"���䰕�(Y�mQ�-�����#|�� �ap�Y�K��!���Pf�;�YJ^u�'��{o6�J]P�(�����ۮ��SO"E�%O�}��K�`�L%큒B��4�+ޓ����S:�\D�_$����S���%��^�������>+�����Y/{õn�&u���Z�+��g,G �1D�f�C������BR��=�"zW�4y�Q���(��`��7bm�Z���/c��5j�c��F���h��#�K�t �
A���*������-s�ݩ��M�s�����-���]���C�.xH)$�"��|0�m= z"�'�{��`p���ń�%��'%�&���@>m���)�GJ�e:��[�w��=WPM��
����n+��!���lҳ���S� ���0.�o�oՀ'V�F �.,�YV �C�A�mT\*��1Q�#ʘ!��Y?����,n�@@���KF��>����V45f�t�ՙ�zT�?G�];�^��7�ZAv��D��h�F��^�X��
[���ԦO2ˠJ�P�P��N^2ۏe��c�o�������ؖ��ثeR��r<xq]$e.��Z:c8踢�7PD�9���ǿ0}s_I�h�iI��������gU��GB�R��.B5+@q�����(��(>����Z��᲌(-��Q^�f��ZW�Gj���Co��	��uPoW\������� �&c�c3��N[�N���BȀk��z�691�Z�8^O�`ZA�<��Q!CB�oy���d��!�D�w��ȧI �8�i�ܡ�?ŋ�#l\B���'n2���d+�n���|�:���D��%b���1 ~$�8�ǥ��qq[ic���>Ɇs�����Y�3�}��N�,8��cw�0M"6�JJ�PC�Q�w����%���׍|�!+)9A�V�IA�Z�3��ru�lD���$m~J�L�w�����^=jN��h=�-q�-�h��K�����Ԋ��&�{��1�^)2�/n�5�;�g;)����tT%X���礌@0ݸ�s)���<� �C��C���iv�`�j��q�L[ی=�J���c����l�Y{�?	x>Sx��]gRY�ߪ;q��h�v��s�'ð�7�^�>��mb,6~x>`��Ͱ���M(�����H��I���yv�Ngߡsu���'@ZH����-0ݕ p|9������.4Ar��i@����(���N�����b��?0�Jc�_���T���?�P0���|}Pg&��N;ޖ��ƻ-���PJ�}�s"�=ɴo��n�Q�.Z�ۑ�;��[�����ba�9�:-G���E^bn�
~\>�_e���sgEo�r�����f�C{,:0�v;��<o�R�R���W�/ݑ�hE��|����B��z�>�[`=<B�;2�n���bňu��."�X�ߖ��
-�Q*���@�54�ٽL�
�Cf!�,���^?�7��?��쪐�����O
F,g��]{��f"[���+�*�rx�
oX�4`|�OώDǌIU���w��ٸ|f�T�����	�2�vZ|�~�>����8�o��K���+�U����J�ޱ(֨���_��a���3QZ϶��m\��Ɨ��<�P��^')ש���rBv�����3�am#�����41�D�̃�C����R���Ս~%[�"�*
ZjX��L�Yʴ���[��x��q�PhU�Ä�/37 9I��!���wf��)��a�*����ۥ��	N~�| am����5,lmr���3WpT޵��a9���,����wV�3�=��:QfX��r��2���֘���3�*��`mS���1��������g�u\g��yP��̄�繼#��S~;-�M�N��1�
,�7�\^��� ��`0��s���
@,1˰�&�!�鍄���%��(MM��h�n B�-`1<�T������P�NK��$sPf�X����0Ŏ5;5C�2+���X�=��AT܃H��pg}���y��G�C�j�BXӂ�wֹ������ғw�U͡�?Z��n�%"�V��e�L��{E���j�c�r*�byc����pi��h�[����6���|���\�7ϔ��K�J�ƙ���_��H�h�����׮��j����,����LV����g���-���	P{m��
��8�HV��J?t5� �ܮ��(`z#�t+�׌0�u+�)��2�9[� �S����b�%3?�I�4$�KNw,�R���NoK`�dR��	��d�>ir����ϔT�����m��I�(Fj�dk$yj��͕M��<w����D�vV�v�	P����x:�/�OUG牳$%���}�؇Gbw���K����P�T�e�q(z�
�(�3Yi?Q�R9{�,U�nG�?YXڬR4��rb[f�	�QB��r�{D^����K(I��Aם��WA#@�ӵw2>��%w�����D,"a_.r4�J�埘��J9A{y(�a�������=9Z�$��Bq�	�as�#G��>C�.c)x�Y��3���4����=��ê�GYi��9V(��=���T&2�K�n�!�b�7�9��׼͞�P`����~��y�T_]e\WR�W����3��o�X�І�{���LI�yU�d����ÕuÒ*�S|�7���F:K�,<Q�jI"��Z,�@���ĥ2�0_l$�:��f>�ftl���n?��j��`�{�u{���"����*;���T�;Z��F� ����1L|>Q2K�Ө�C�x��$��́ԑ(�§@�鋦��U|Ր0�SKXo�K�ѷ.!2"�ݶ��K����R��%Y`�;�J�L	�% k�� ���p�QY.�������`�<��#-4 ΐ�A��	5uڿT��`J�s��G��N�	�ȱT}3,�."N���M- �+��F$�����f'=������d�����0b�h-y�9����G��F�-��n�2H8�@%1(�Ft�GO�7wZ�](D������b8���9θ���_}q�<?��b�a�~�� �Gߜ���3,����0q7�쟋��k��#jnb]��`Â����8!�Y��D��G���BA%���f�+�o;oUE�Ǐ����|ny�����q� �	����7����ä�j��H�c��AFj�������ˠ�`��ܧwu�nKn%+���E�� �.o� 8�:S ���mu@Wu��Z\�� ����[tSd{��Z�h��e�u;v��K�A��v��Z�h3}�EJcV��.#!SK��?^����Z�І'�h6LcE�W���E�D<3��H{���m@��&1K�{)0�a_i։	���v�hsʷM���1���U�\�?9�P��[��A�P2������n�����@�nx�T	��,�� ��W����=�Ag�B�ϔ1�m�'�~�;���d�;|�������&c���}O��7c�T�P
6�G�L�
��-�#<��LE�A�w����U��"�[�j]�
}*3gu^�	k��$X͠>�
H ��]<>�NDe��Ӽ���*�!��Y�!1��f�i=�ӸoIfOz�#�?�2 �ծ5�?��T:��=sϫ��`Gq�5�ݑ4d��i?�ɪ�7Y��̥��W�AX��.��SO�d�BAh�7R��&5���t�d*o����!�h"z���$��i�=��d���wH���_ �f�{#tc��'B'�o�c�ݕ�~N���5~�Ǐ��7���;����ZŁ�o��UE� <��[�W�C�!f&_���2V�y�o��F,�Nv���e�d����*�bfZ�Qf3��t�<�$��,����}��v@.��,5��!=_=s��M�����ٯ� �ĳ8�l
#��5� �F���x��oR�N��x֚ ;3�>:Ir��`<�I�V��J�1'�Z(q$^�<Xe4:*�X��D�x���RI_(�u1P��zG��֙m;�M���gD�Ƥ�fMv{9�S�;Z�vt�Pک���v�����Z����^��?��s�D�T���s}�|���p�4`�1ͮ̚�a n��t�?�m�o��m�,{ ;�y�������^��g�[5�2'7eB���
��&#� �Cr��3�Te�z�һn�JM�HL,�Zi��oi�ޫ�Z�;7"K�Lq%h����?$oi��2�U_�ܠ> ���с,�7<���hp(�MR�縮sN�Bh=.9 ���`4�7�n������aP)��R�*����n��'kӿʬ�"���(i�b�Yzĳ�\����%�	5K�VP�~�d�<b眺}s%���Dzf�ElptQ	`�X'pA����%-԰�G@��ЀRw#�s�ѵ�M@�R��b�^Q��/�h	���	�"�^eR��>�@N��H�ģ��i���|u Gr�P�i�wH�.��tU�ɷ�B�Guk�n�>��H�R��~��G����������ͅ3�����C��<}՗~B�>[|+:ҔX5��q�` o��%�Ҁxl�Vu��m�����l0Աrm��O}Sq���_st���B�u�|�#Q8
j�x0` r-�v�� ��Meh��`���t��>�7"7oZ ��
CY��Q����\h��a�濄ᒚ|�I���-gHY��~��/}ɡZ�9�4C��EP���!JъW���"2��S\S20���冺h�)�;F?2c�]��%��,lzQ+Uu�%rĲ���j�6<���>Ў��8���Ҧ�m����N)�b� �\�f�]�+�v�k1$�w΁ov	 [z�v{X{㫊��r�3�".�Y���8j�U�'���2Ea⤶^0�pk��K����v��z�B�[ ��%XT�Qk� �w�Fn���d5�W��R}:���&Qd�x"nF��-��2#Sl��Y�Y�$=�a`�,�-���yE�5K��G�hɼ��Sa/��*6� B�<�dV�οSl|\c�����{K,���(	��e��ٱ�0۽$�yD��~i���K�\3_�����kF�mlL�H7:m��98�����=��_�������y���9�����䑃%�**���P�W�gI�p>"��'�FՑߩye"�G�&�N�~�3:�G�~�C *��$�rRĬ;�|q
c|�A��	(+7�>1�}+qyy� Γm����A�gP�,Eq
j��O�tcD
T=���)����9kmh|�T[�k��a�f�	�0O���6,����(�n��q�r�'���tٙ���~iZ�z"�����Cq�ٌaUt�����}�)�*�!�	OF~ĩ3��1J2�6��-鼩9oX���0�D�����9_�W�њ+o��t z�}�
?~�``N ����b�@�b)�zV�Z�ڝ�
��g-n:\��Nl�����J���ۯHW{��yYV���%3|6�v���������Z�UQ]��p�'	�Pا�b����Cm: ���S��ɝ��pD�=������r+6�؛�����E����M�	Xs��]�QGo�xS�7Ი.����*.z�h�Yh�F�tOJq_���ū8��}�@A�4l�Ic4��8�F��V�ָ��5�n�wX�A�{y�r�F�tn��^VwS���l.��4^��bI��d�҈�	s�_�ٔ����J;��[�7�����.�͉��}ۜ&��S�W�+��	¸E����|,���jk�>��o�z�}h! ��2R��`�,���a�l$��I�(|fHڷj_��P0�[㈞�����F�{�������K�<�+4_Ӿ`���\%��wO���QP~R��	-��Z��l�CUY��Q����?��{>.兪������qp���i.��Zy��.��X�f�cK5U�,�fz6���+�Ő�u/��L�/啗cɕշ��y�hs���l�@"1�E�R�i���c��|��l�*�V!0��!Uغ����G�>:U�m�x����F�=�$��Al��7o+GnD�V7� ��:8�� 
;���A'��?R�rit���hk)Ǭ7زnr�1�{Y��UXxyxj����*,m�H�W�Ioˀ��>�S�0+�����2���t�af�\��2,�}�� !�w�P���~�Z�3O�	sGi?3��v ����I���j��ATl��4��A��Sq������@P��>d]���E*2�E��h���<Ф;����2���\#�e� 0� .$9iC�c�ϲ��o��=F-%U��ZIz����(uaΌZ�%;N���J��t)��,ah$�2ɕ��iOT�f�����cr����^��M3l#�'��~i��Ǌ���^xx�75p���M����z�jM�<��`��%n`]�>#��q�3�Qc���\64�M=�,��#?UOz��&/'w�{�ڀ�o;)
��eI���ZŨQ�x���ҩ�9{�k�[⸗��=�������7��^���f;�}��D��{cx����x����B�G��D�qeH����3s��.,è)6X�w9y�?`�o�S'h��͉g���O�p"�A�9�"�0c¢�����B�Hau��G��&���A��"��4�XJ�0�c��J�d�i�V����)$�Mj\���n�>����?�7��}���\/���vX��H`1n*�c9#�_{���X_�u����V~T@v٢��4լo�=����T,�+�����h9t�0���Tv:�l^����zQ�mq��@?j�e�|,"���e7�ΰsn��XL�m	Q���Θ=6��m��{�_ʫ!qg-��^�,k*u�V��2��Ҝ��>Rd�*~T�� �N�"���-����:���Q8͌�c�ӕ��V�[_4< 
�boRsijg�46ύ�g<�ˇ���f .��Z��U����~��zi(y��P�"�	9i_� ����Bo��$t'�]��yG9�9���z��1��x����+Īuc�F�E�e	�EX���(�&p1ށ��	�򍮩�H�F�g�<���g�Z�@m���@GV��l�� �S�D~o������29�U"gR�x�b��":�ǩif�5��`��J.�ݸ�2�q��5���	['Du�*-f����//T����B��
~	H<@T?��� �c�����9�:	x�ER���؂>����f(4|�`<����<�^,�I�d$�"�=K������:��E�4��c:{ND�u�#>�O�Z�G���g��h���)�~+�J�#t,�c��8&�(-a�n�G�ŏ%V��y�D��e�ӆ�:U������?R;�\=�-������AL���d�m��t�㡁`�ʹ��	��1?��<��EV�T�9�1úGtT�TJ��K���~��*{��˛��ر0���	[ eR��$���dݝ�aDZS�I��L2^�v��qU�a}�P3V'�?�����橭�^�@Dj1@���Z��ݥi�\7�B�ڋ���!:���@ǰUeW�a�rO��=[*5��@����:\��7�R^J��~�N4�6ގ�8̃�VRg��.��4uN������c���ó��\&���}�f��	Y�
��<^�8тU��p'���*�u^��}�牙4yq�����4��W��݀�����a���/vQA�;�����_~'.�� 1_͢n�����w�4��J{\a�kK#J����0��{�����o��C#)\${���Q�7�6�X�%�kϴL��f����{X�3\�ɨH:v"i��3܅5��#[�Hj-����~>��m�	���Ӽj�l�˷�!+K�xJ9�K#�L��̋�qW%p�(�U1���B�Hh�������z����7]gH��:'�v���nFIOY|�& �y�R����K�7�j��dn��(X��:}9M��.͗�0Ϛ��Q�i�8� �Cg����P�G�hT����l� ��b�U��}l@�[Qf>򁔩�A���`�p���)��C�ήC	�A&�B�ϝl����f�mD��4�_2�D�u'��/�<���Sr�6��%\���^K�Wq~S�PH�b�v>����r�&Bfc��<��"�؎��,�� ��V����X�lO�}�ݤy�?��%��B��P�cF��@��]7�L���cHܔ�	5��lE��v�g���?9���������6�Fg�p� ��
fK�KxÉ�6��!J���-W��@�3̃��Dɏ����� ,��@>�@�O	�M�L:��cԭt�
s��2����I�Qt4�d��7�u
O㤥;�4M_w5j\{�Wy!������Op�C~x��`z2�����;+�s5)g�ؗ�,;,_�D�ʊٖ|�F L�3*z]~�ꇮ\����#�W�&����� w��Q0ܟ3:�=��T��r`����o"X�G�k��$�L������4��ͪ"�wj��F:�8�Ok�Ե~&�ybk�m�k!������&���^+p����1�:��� �z`ފQ��>hqt���
��{c#()�AN=7U��$i�;̝�}Q�HGW��U3�Ɏ\s�=��V���rn�+�?��"DF��5�z�M����i�<�
�ےz�JB�{�T�9R�La�NP(����n�}�f zTҕuMK18�)�i��Fn�R1��I���|$~i�Ý� ��,�iN��&M�V��ӊ��0�#Z��b?իC�75]�����kԏ���
K�zn��	ȥ��zL�}�9sY�w�9��j�cR�=����$��ɨ�x�4��t/�5�@ȳ	��J�u������$���bCb�gݤa������G`��w�#��%�߰�5'�_~�E��gٟ8V��&5!�l|�t�t��(h�ɏ��������u�������G<��;��>S�����x�q���&A}bj�(+�^\�7��M�����W��/�F�覭����O��O���&�2eI@-�
,D8ΖE6�3��)�l{*i����[��l�Ox�;(��mr�P���W�H�-������Bn�w�O�ln/���嶝���w�e�{bBt�+�(��+ǩ�~/���
�{V�K]������ON���cت���l,)H�o�U�6޼a[ׂ2�=��DV?7�v�Z��Y�[��F��9�Sq�4�E�n��$ȼf4dH΃�b(�N���������M�z���¨���p��s�4J	N���bb;��S��D��Q׍�8TZ�&���8"�����{�3�a2s<��1�lJ����0Cx���8��4l����:Q]����9@O�;��0���%1�'�j�y�����;�~�m���Q�zc�| ����J��|6R�!D9��J�o��kR�o��s5n�(���ilM��/BAzB��:�L:|I�D/��чN}3>+Z��}���������K�,�N��h����miI8�X�@A�)߹p�k������|T�30��#0��HJU�=�6 �fQ[����4,�?���ক�JsZ8I 0�\]���b��z����ɹT��*v�	�޳�h>�(��kc��	���5Ӗ(��m��KS��}Q�ABo���1sOO�j��h%�j[���%W6]���~h�u�w�Rc�H�z0�ҙ��}L�V�>��xt#Ҷ��ͽfK����Yt	,�3���9���jݝX�s>'�����z����3q#��h^�v��9]1�sBy�Ѱ���m�d��^�Ӄ�_	*ͅ%��l	z��q�\i��!�1��hN�d���4���zy%G�`P	��R�hЬ�Y��5�~��Ţ𮰵�Ȋ)��j�����X|�P�0Ud�5MC5<��p�@Q���c��[76K��%6���'|g���ʖ��
>���E	��^Y��Pv��UѶ���"r[����E7�M��<�ɒ�K�%�5)X���(<�t�Z���\�f�U�>�̤�F[�pժy��JQ�<�Q�6�?�|Eoh�;[��.�!�3	4�{���a�_V�7�o�e�|�a�'7C��r$Sÿ����|�/� _G����:�wc�o�D����T�R���N�`-~Di�^��\���0�3�y�to�M�+��D}1�G4�I���!�>�T�&�	9H�*��~��g�Ӯ&aԞ����p���N���H��������`ao�T��=�����W�BW��r��~��:�K��n&Ț ��"�Z��dW�6�m ���㕭� �#�^i2��a���N��p/K�V���F��F�P���g�9�fO�tf$��9��N�ϑ�W ����"�͍�_P�����ԗ��K5�y����\�~H��jW �)����v��hSP��ʣғ��B�t_�K2��G}V!����4���MҺEt��*�HkH�Ym/�ғ|87_�Q�Q�s`(��Uu������������n�Ջ0��X��S������D���>'�~�1,zHgyp�����|�Z�r̯� Ũ?��#E>�J� ��p�cw�\����p�^��fr��<��������Ore`H)T�Q=�$L�تQ+����G�|�K̕��[ �ڝi�b)�ԝ#}���Q~nK_�d\[����G�*Ha��hFj)+���k�x��䕽樅�MG'�Y��Q�����֬
d-;�L+��JZɶܤ�ԱH>������Z���\����g{�Q#��;��mՐ�Y��_�А�~dfR��bCo�?����L��&��bcb��g�յ�Q��UO�f����]1%jmC��q� �#��;�.�Bj��h�jW|���X<δvQB��md��v�h�tFos����Ta3<Z�<����8S�����G�8�n���8J��il$�eu��L9ʰ�K�6Eh�hPb���j�cZ���'��>�f�d����B:�'����QZ���=��	q�<dz�"=w�B�B�gs��u�t�T 1O}k~@="���*���#�Sў�L�y�Ys+Z� �c���P��ضE��\�l�t����5�eo�4���u��k�K�,c�C���R#OO�Y`�d��X|�1��{�;�#�Bl_]�[ Db��xE�e9�bG�j��S�3��b��*o�8#�lD��U���:����U!��n5Fᆷꢷ۽)�!_!����օ� �|��`<Y4��^��	�D��(*:� "��:m��K���Cō\Q�M�;ه�q)�X5�qc!'6���Z���_rZ�J.�l|}���۵� ���>�Fk����Ia 싖�� [:M&�jY~'�|���r^o8'(��*�|�n���9HW+r�	�������f���y,}��<)7�Ǣ�r�O�]�h�X+� �Ɂl;n��k�<ױ�'v�*�ZT=�����@WT��rF�4����Vm��*d~6@����;���4������LP���:�V���
�2���c�[��S��k�]���\I�s�R8�u> !���:�S���ec��]�q�o��U��%9"��B�=Ã������SC4A��ا�X\O����+�7��{ce�a�ל�ˎ��j�.����B]s�A���~�Yt�Q�O3}Y�J�J�#;i7��e�irʋ��E�1&[G��b�Cg>�.P�[?g\�KKG�k��@3t`��<F� J�ev�(ho�NY軎.�!h�s�� ��Qb��� lRlo_����#f��(i�}Cn�]���0k�q���ɝ��7�+�br�Q�VC��`܍��YO��͜��͹�@��H�|�& ��&v�t�c�#%Ez�qG�ݟ���llm�w�~-�8�U2�v�ҋ�.�K��CYG��k��w�0�m7��h�t�2H�r�z���ސ�����r��g�v��eM
X�EE�f��¢�_����J3F�@$y��9�&v��S��U�k�S��\CM�3iq�g�U���nқ�-��=��}��mÿ���DFLG����T�{�E{ҕA�Vf���k���q��uE��E�}���_n�ZEWY6Q��`��7e��/K|�O�V1�XGr\���e����o�OZ��J����Cё�J���K��(�2ګ~<�[��h�\���C
�ƈ��X�ĉ*h^��J�X���N�wr�W�?��O�%��זn{c���ְ�=߀7(��\��-N���w�`�O�ڶ�'�)�U�]7�N~!��'u��W,�h�F�ͣ�'�J�q��Yu����.҅�)����"03��,������96���q��⊳<��,���
�׈.�jl�&�>�/*�����v��0F��=�	7��
����CV����J�`�<�1�q�������V�4��(�K��h��!ɓ�@v�S��n�A+j/.��[x�MC��=���C���Z��,I�� �8�cI�n���.���V^��(H}�	/F�R�˭��C·n��ă�c��i��<�	����% G(�l�.��d?@���L3|��P��
WA���J�7����po���XI�!4�b_\k[�8��Ĵ/��So���˪��A�	OU}��,��
�OIvT��.rw�-4w^wv����ż�ct�/��s��4�D�����E����}����+�@~�g���N: �g��*��1��
�C-7cA��d�	�z5�A��M�2v��l������>��S\R�aꥸ"�|!�����:�ڠl��� �w9Ѹ�]t���L���łJ�6���VWΘGB�B��a��ӯz�C67�r�7�l^�z�G��)�^.�9�E�.�Waܦ�����宇�0�2��K�Ncv4Q+�E��T~Y�On%I��OQ���|X�T:]��%+��Ap.FN���ύD��_��mwdX|!�O���R8�C@�PQ�ɵD��
��њ?kY�m���(�;��m?r+u*���|N����}i3�w3H%q��4�C=S�z���Gp�<&�[og/���6�%����@Ieg/Ȏ�ZLZoԄg5A�c+�Χ��XF��}� ���ɮJ�鮤읯�1�6���z�N�>*V3��n�7�|�B�>����X�)>KL��֑������$�Ō���2Y�K��� �FߝS5Ux�IB�g|U�����7�7g��Ѹj$�M��\+�O&�l���#!71c0s/WK��Q�����? �k�<	?
��:�@꯻�f��kg	���pM�K3�V}U�V�����a�����[t�[T�Y�M6�*Z1w�&��EKn%a&=��ʹ��}J�ĳ$FT|'�/	F"���(w�R�˫��I��g� ���i[`��~D{6TX;˖Sٽ��@��{P1�B�=G)t������_��F�t�a02���ǚ�6����)�W^��f����H��{�y_��3&G�ԑ�K>+�9�Ԧ�S�Yv�5C;�sX�`�3�Y!,Y�͎S���ݢ���<�/7F3��[�� �x��C?�U~�	Ib�l��:I��5��I0�m<��[^5�H��G%@�V����y����L
�w��B�5�d֩1�rx��GZ��	!��s����1�ថ��p��Z�k?���x�	�g�j�����:�xTխ�$�Ξ���S�	M���#Y�����)I���K	؋ڤ���-�~�YsXk"���Ԫ��D:"�wIg�~� �Tx?^�j)2�.���E}i�W@��)�ϵ���|)V]�C�	�On�
���E�����nP��h�A�6��4�%�[�ǖ��SFa�ur�L�M��U0���Z�0SA��a=�^�O���	�F�]Rř����	�^-2��E�E�=��i(�!EEjP}��_;�eU�B�����Z��xw8�kd�I�񍍘���1T3PL�v��NS55 �Na��5�\�d)�����^S&xgQ�`L
��Į�}����p��)�;�@��>�/}޶`�HU��NW�c;>��$m`t���g�_Z,�%X3�*wl���UXh#����[���?W�)q�8øx�;i�H�{�qn��B?l�U}�_�G����7ٛ;��Pp�n;u���tD^�~j\'�(�T*p����4nj��V����ve��c>����B]�P
hG�o��`�֪@�Ԗ���/J�mt��*�v�D^N�\��y��	bŖs4�(!F8������>��VƠ����
a�ěc��g��:2���PU[���25����<]^�ڧvGFS���Zɹ㺀^u6$jy��6F���u�)Y��c���A!� ��\N���T���W7� ���Na?�I��
^�'`i��"NTb5��WJ�Eg�|�m%3Ƈ����l=P�R��* �j3�����W2����;~�=ߪ�00
��J��5�s�#�w�(ȴ����˶�-� D^*\ת2��%�A������Y�kO2u#UVN��rװz��K��`���W60e�Yk����
(�ɼ"�=g'G����o���(�*r�#�������"���	�q��߹�U�z,Vs��I�S�^v�T@�;�f��hbw��� ���Z�t	���`��E)���[OjH�&�g7����P_I�O��� ����嫭-�|�� ٮ+D�����>��ʣQ=E]�P��kr�sV��v��St�b�9�2sF���8����/r(M�~F�b"k��f����)�:����*��(cO�L�J�;�
-�e�E�����41��f�X�U�uK9wp�.�R���B'�&ܼ�˨N%L�ƀH�Z?��R�E�cR��dղz�����Qe��=�q��،�Զ�SE�7�K&��r6E��}�4cJ@2�D�+JMIj@���M߃$�*e���"���3ۻI�%���5:�>��H��ꁉ��\B9�C¨9��:��!*��o� ˈ�걃���m4���-��*�2���{$/�F�|,����k�])�l�:	q��îR� ��Lob���f�K�H\��l����?�a��t!�@�Y�B#�ٜ�I[&�����d���z���lKylP t�M�	�~?T�.>�ǳ��?ys׿��j����k�~�/���W�(#W���<��]�c�i��<1@h��	J����=���3��åw��ѽyn�;Jk�
��ậ�:ɞ���ӬX'7Ok[����y��&����Lm,xJD��}�����I/Z��Մ�˃%���旇,aW2��G�O�I>��b��η9��9S���ί���!��c���c;\q��l������G��q�ؑ�Ǿ9��]� 栀<9'�P�:�=���l��p��Vz
:��'��F�V�]�ݤ�K���v&s�7	 m�w@�ki;�!�D5j��;y_Ե����V�s�R]d��*�p�#��1 S
�r���Wc�n�|��q��(�]gF��T)����D�>%Q��J�$�&S�Y;������l���Z�N5�L�@���L��[�#*ு�.��"�BiG�2!L���d�N4tY⌋<��z[Z����I"������;h�� o��kw0�A�ޱ�[����^�T�_�!�lZj"�&I��Q'WA2�;A�냸��i���AN4Z��8*(��,3v~����`k����DFg�>��z�xֽ�ouUl�q�P�*���
�:����w�����by���bE���S�x��⊐���� ��]��Њ�!�� ���gJ�HiB�e����-gȦ�c�Y�,60��Uf�E��K�ҽ�d�G�=��-�wà�/Zeιa���	�q�P��<d�<�	t��b� �c���!��{��X�]�4���I/Ҿ�]Pi���Khs�'�����¬��@?s==	KK��p{��F޲�#L��Ok,�*G�$
`NO���6��H�_���Y�f��g�iGԉ@�(斢�7, �?H��8LȄ��ڊ�����i� ��Ʌ}8�V�}�Ͻ���>V"^G��y8Ӌ�z�P/���4=�n�x�U|�7RclG/��cI��;+��]r���!�jJ�Y[y��`���+/��pk�k�V�-%Q�N�9�w��l����G�k��]���}`���sT���	��G�d��j*�R7���� 5Z�۷��ɵɧ���8�L���F��X�V@����j�˪���I�G���8�_�����A�ʮ����j�M����\���ǧ_��k�B�#�j���r��i\�:֡LX�r6t�n����bXp�wg����)�_Zuǎb����@�N���E��{��~a�y:;���+c/]�7Y,�Ѧ1{r�:��>Cx�� ��!�����#����R�k*�-����k�z4٭���l��f�~��C�yUN�J��I~�?��#C���oa��I�"����y9)ͳ��̊��C(+3yq,\�2^'&߱l�X8(��sӐ�%�I k��A�_��n��o�����<_l8u�c��<�1 1��Vm���LB.�n �1��
tw8�zp��$H�Y��"�I�4n���T�����7�U|`����q��W<W���H��a�>ֈ�s�����D�!��9kN��X&@!l��x��+j9��z�8����9��/��&�a� �̌����љr�5�@�Y�W�Ѿ�Cv�ԭ0?$�7�^w�<e\����m������C-B��:^'^xd0�����qz��lM���(tF�N�t^I��-/�E+	@]��,]�VU��
����ֿ�Z=���G��t�a�W�#�{�����UB�%@@����z����щ�K�\E��*�g�P�Ҕ;��q�M��7e���X���-�&Ȗ�w?E�{k��d�A�k�z-���$l�������0�ᰴ?�b��d{Z����gJ:U�_叾��P(/���!i���>]�^��� b����]ɇ�m�e}+m��[�VÁz���#�cpA��}�������b���,Ö��#6��/����~`2���M�LY"H�reCF����%������$�:���R<�\;���׌p����N��� {oQ��Ϗ��x�X�;H��C��ځ�S	�	wC^�ӴbA��g9I4t���y7.�#�`X�݄�ԍ6���z��N7ɩ��A���%u��*~�������V�LH;�m�' a�)	^���$D2Q�R���>L,�V��Y#���I�Ә�۷�z�6+-�"
""T����de5ˁ yЅԉ�mt�K�(��S�9�N�(BWd˦��*��?���T�@f�^�d�l!C^���i�O����S��
x��%B�[Z��f"���8�G�O����ҏ{S����㹁ynw���E:��:H�)/z��c�z�c� 1�jj�?���"�d���ňTJ�>6��H�ce��L^4]	���m��l��R��g��F��It z
������a"�s=C�h$�/���E�����!'�z��Ӫ��`qz��E]�\� R�q�IӐ��po1�),��bs�Z!$�	�w��`L�<�#�)��Q�ƔK�aa:�9f�9� O���+_a�lE;��'�_���	b,��k�s�Ͽ �e9���S�
���5p(�����w��td���8�O1�	��u�ڎd�U�Ѐ�&2t����\��°u-�a����ݵ�r�ma���2�r�8�V�i0�Wo��sunof��-�S����-�Z*�0|x���r��|�I/�Rå5l}��
�l�S�Zؗ��kݨ}pyI��[�5�xG�ڢ��:+3�b�����	��#L`74?(�K[}�ԋ`w���'�s=̦z���y�>Tׁ�H�ą��iH�:/��~��_�݊���N��S�b�A�>^�2���x��1���^��\��hh=���� >6�D�
�����l�j����:�˗�;cN�/
�E�GʜN�;�ߊ:��=\�^q���|<qX+)w�w�Ơ�)�2�5b�\����F�X�����߈1����������~�����#N��W������SD2��,8ލ��m6{�c�R-U��4���soۡM�ݺ�$�
��>�(9%� �\<��U��[��e��z��a�s�!W!Rۉ�{qؒkI;�"�Q�h�k`����M �M���7r�%�m�87�i�q��R�̎h�۟*�/tf���N��G�(����Ta���tB��ߎ���&�����?����d�w�������
	i;/�M>=c�F!˟vX�Q���Ō�[���0�;![�s�;�	�j�׈��p�&��w��K�}G������L�������+G�rg�+(��~�ף��o�̱�oL�oiGd_�L"ɖ؄��K�YAi@b�<>�t\⚵+s�:�	�ԭ�߇���h�O�$yzaKr�z-�!�Ms�V��/1�8��i<먷
]^�*�����K��'֏�ï9��U�������N��f�r�y �_N�����%�=���������v3Kڐ�1dj���C�EY�g�U���[��;V��5[�=ޫ�_��㓵
��|��)~{Q�A��m��S��UUrʳ.8�hO�R�_4��+���J���Cd��������J6�Ե��骟��	��n�#��Tw�O��%(������R���y�*��C�	���ݥ�Gz�����L��r���j{˜�ྯ�r 3FÆo����맾���ɝg�ċܯ�k_ˀj@�Z,�QUS�+��FNZ�*���HO]JZ����I�*��5b�q)!�+|�����#C׾Dl3�O�Y�V�=$@m��3�0Â����� ��e�>�W��G�Od��v�y��n������s� 3�9�UQǭ�Ơ<bWჷ�O�f�^.K��7�'>���o󋳽�*�d�yƍ�O����;�Ȅ�F?�O���;������ǔ֯�jSOR������ ��Q+�>p_C.l��1Dx���M"?�¾Lq�2PZ4E�����^���}�qo)��zc�Y
��������*2�hzxf>hi��`I�S�[��bI�W�! Fz��a��
��5b7�5���F�dD;��!�ä��J�ߨ���=b/V}�zf�y'�s�*rE��>���_D�IR0Bkx�u}�y-�$+�������O��U��k4���#A�M���Y/�'�1�7���N��DJ�IF��7�}i1=��%���f�����%��`Y�s�y����駦�B�9A%��ˆ'������^R���SP1��Y��QAi����ق�����c3�'��+�Bٲ��Vk(S0%�u�6r�Gl��E�)}��pB�h�J�Y;�	>�^�Ͳdx=F�X�Ӣ8�U�<h���3��S �o`p�A�n`S�l�/�����;�vp�>nl�z
�d��O���Ta�2�K#�\ʭ���6�\E�����k��!0��C�~]�C�յ��� F.�@����A8⧶�Rb����rpl�`x�4��-������!��vU�&�(>Y�{�7�����cG��� �~HrF'���������8�4���7�Ӌ��zy�Џ� )����)i�� 7zc�<9�AN��8S�1�\eoA�J�P������>e�]D9]g�.h�C��Ǔf�h�O��|����}�M��뷻����ܰ�ni�j,���g�V<m����'	~b\$`�=dL�kF�п�Y�����U
4$/� ���Ձa���^�<�����d�u�-�Ka�|��jDJ��9�[���G1nb�P_/ez�1k������Y���v7U&�%�A����ǎ�2���2�'��Y!���*���ּߛ���,�B;� =�B�?UR	@��̏���T�����d�潕��[��ჰ%��%�u�Sy-��Xݟ ��s�B��[����;t]��9��ٗ0�m��R�ɖ3�[���W�N�5o��A��10���b�����]�X[�H�i��։�.�:��3\�W7Vlݨʋ}����V��]$�BYIHE�T��Z;ȃ�=	�K�98*������C^�dX���et�ʎ8dU����<�d��I��}:�Ӄ�/�5����0��+����`�'pZ=He>;�]�k/E���ϛ3�
���ϵ/�xֳ;�")m��sw
�E�p#	D���_�iv�
�M��]���T�a
\:�Hl�b��+�#)F4�*m�Z��o/��y���-P\
�)����@Т]�'�zn��"��j�7�5k��}l��v�px�;��k�#�L�]�J�g�ө�Q��z�jH>TG������$i��uh���Zl�Z~�4�цd�Da/Q��Kv�*�^�L�z\�є#=�߃�"v���u^Y��Ӏ�~P���m�;��x�p!e����A]b}��Ѥs�r�'R.�8vXZ9�X����������Hv$��ؕ��9s���7%?.�_�:���P,��^�"��b�7\�