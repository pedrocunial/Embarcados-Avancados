��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c���ѢǓ2�Su���;���L�X������8��5~�������k�Vk�T�%��т烰�{�r1�������E!� ĲB�Y�l̮��U$�Rn/z/G�kh_�id� �i�["���$�u���%Y�@���ݨ��DxQ	!�"/��i|]Ag���n�+�]�^4�	I#�P�n
V	��+p�զ�~ŷ]��n�d�����>8�Q_Aاc��pgw��!�ǂ\e$f�v_p�@��G(Tf]`�W�,w�Yz_O&�A��
+��C�?ĉ�zz(���?��:�vl��g�qv��#~�\}�yR���*��vmh�I9h�*�/����ǖ1;$��a�����N+	ݥ�.}b�v�2���M���QŊ�{�"�7�pmGH�˃-B�����;��*fģ<;ƼgX��qN�����5�£�ӳQȕ����IK4��̣Oc�fQܑ��=,5�P�ǩ�}V���s��zބ!Iɚ��ߕ���C/z6��in�������D���^#J�9*�}�N	�� �i׸yՍ�:�D70k-�.�����jc_îA��$c����i��y�չ��?��q	��_(����N�몒QL�^�mo��ĀP"b�@-�����^F]��;�ʃ.3E��}5��9�E�h)K�&��j��!��j	g/��ȍ�i��������z
�D�m��/R�����:;���C)��c�n}v�={��'w^ȿ��To)a��
��'Y��{���%��ɺ�]��O�5C$�~[��o^���Zm=A~���A�"Č"*D�o��ecQ���{��HQ�؜��Fj #|�[������l�3�ոX����X��%G]�fҾ3�:(}bU�޶�E����D�:����ͽ'ͻ�g|y�d���K���ߠ���jL� 1�-nRe���w��$�y"qa�M!G�^����t+T�Äv�sU���V��ʪ
�v�%^F����B��=���.C=��msLG�2� nyi�-W-	�T诞D��q4Qv��f��Q)���c�o �%ϵ�<��!X�85e)�=>~�#��d��%	��%i�`u����c��!<��<6�ՏVM"1�}����W��m���Xt��N&3��r{S:^�O��H��=���)��
)%�������ס�5ڋ1���;Hu+k��Ɉ��W�)�ͦO������8,xQ�*a9%e��f�[�K���"�x��
����K�q˵�^��l�F�I�Mn�(U�9�g^I�p��B$�v�m��}��{7��Ʊ//��08E[�aG,'���ke��l��@���i��֞�z���`��c3.��C�#��馚ŵ�R	�gI���a�Pjz�)�O/b�+#��a��hA�����\�p�P�#��8��j�4�mq�=��N��_�}���$[�U���� x�����b0~��	b?x�B��e
x�>,���kt',1��������q��B~��r��k~!w��K�'�Ϧ�T��,���hǘZ��?���Ǣ&�3fF�LB~Ů�Vw<��s��ū�{H�Cyá�:�n�`���!�F��$��Ka��J=�1{�.��;1�O�ΐ�sL�d�W�ŝ-89,��nuCac{V�E]P�8}b�A=�e��@/~�l��ȉ[��x����?J����'ޱ��5<=ܺ^�hG��M��K�o��)��aN�h�7!��5�I]�ɮ�4Z��E�+#�����ݙ~���2�UҸ#��[[���5}�By���Ʊ�2+���K�g��-X�%2�F�)�����U��`_��� c���}�|�6��g^m����L_v&��lgji ��	�,��Xʀ}4wYFG	��`=���P�lIYm�ve�<��&�H�\k
6�l}2W@Q7)��E�47�$m�?}{]�o߽��%�p�E�Oe�� �%L��m_�z�o�������T9�q��X�7����U;-���(b��h��Z��5���Whm���#|K����=ׁN�I(4���^��%�0�yc�	pmT}>I$���o�)��$�"���Q��O����e�v"^0��T�x�͢����81�۵��桞��3\�{B�xY���s�#LK���S���5B����6�V�Z/�DAm�+�im��}Q���n̷�z��D_���PXɳ���8/@�� ���d����Ǖd9�r26Cg`����k-G*�|cc$c&+��0d�5�^)��83�4��K2̄�.�*�wKn���Ѧ)�)T�މ�-oQ�tƏ2�_?x|�= ;�I�������A�K�g������-=��~�7W4dh�v�D�g� ��n���WE���Cu����s����Di|����+73������c��нG;������4R,|ik�cr�+J������,�����/x,����|�x/_Gb&�j"H��,�I��;�"�lP����F�H��9�{�g�m,�+ga՛S�fˬ�=�mD�O���OX�u @�|k�����r��s�F������Ì9���9!$�M'#�}�%1�5»GiEen�Z���
>�t�������	���!4(��';�y��z���D����I|� Ϊd'��׽1L�c�[�-�p��:v��j1��_&��ޝ��}���O���o��W8�0{P2�5	\�8�޲���k��Pi�y��C!�u5Y+�{ۼ��B��X��gB:jJ2��ep�gv\4kұ������Nx�~��h��Gq�V�M��6�]*X����x�L*B�4���֒W��`���!�t5 M	Y`��|�����>�ʈ�n���x�Ԟd���:�hV��
��J��z�
�{��|ɱ�'|���J�[Bc��\�`��q���_/��Q\�q�S�rf�yj�G���p�a����!۝��ժ���8�*��4��	�@���?�����юz�&�	��w�x�&-6�t嚄*�3�moR{Z�`E�P-!
�x^|��X�5l�)�
��xD�i@m�Zl��t��gn�愙�I��gS.��wN�mU;������op�kS�� ���5�v2ӯ"��i���҃�`�eNi���q�B�l��-V�H.���]���~ŝ���W �\���^���{����W���ͺq�<ͻm��.y��!V2(�$}��3��|���	���5ةzN#�mᢂ;��2�"���y�vku[X�[��o$���-ҟ[�e��z�(-2F5���Ձ���+���k�C��Z@^74�WmA�RkG3�
㨑Z����v��F��HE2>�8TKG/�Q�NOu�!b�
���vq�5�c��O���y�o�-�n�m���Oq6	�?��^�ߥV�V+;�
��'͈|?�D��P|�y�T@�wD�f�8x@Yj>�0��������A
u5�_��n��ar3�">shD������,�e���6j' �$m��Hl�����J�������I�$�p�;��_ ����ʟ�I	/�멫�OP1�c��"�E��$B
?�87s�Z;���rm�OF�7s�1��.*$2�u/i}�7EðH��NEv��)Q%-��f����@��P�.�t�Pp�Ц�o��,���+�9(P�޾1�t԰��3{B���b,��8Y%ʽ��`�������h�%W}e:���f��[�P�p��I7�:sV���? "�n?]y��R�n�\,t�k��S�s�aL,��E�B���}�������Qrӑ��0*��a.�� ��	%�k��shT`�q��19_�%�zu�3�i�ߺ8�/���Sd)�Ӻr?Y��~��U�|\i��&�͢��T���x�>��?7T@��r�T>fڴ0w�%c�0!b11�$+ŲO�E݀P��
ْ����\��/Մ���l~
���٤�2�P�K�+6P�,>Q�M���{P#�ݍj� ;)'�+��mO�v�<���O;��(��,@�	pcm���Ēf�D;ՋrTO*��\�Xܿ�ؘ�ͻE^��E�(�Ao[}��
�������ZL�\B� �v����i1� ۟ �72��(е�u ���Ny�?ό�3���{�D�Y�&��vd��*[5�f�m��4�7'74��ilu"6�tn��M��nf���kA7�����9�}���n���[�/	wK�@rxS.YG�s{�A�"������]�[��bw�����=u��¤�1;��?�Tj�x!B�<�c�	夈��iՙL��R��m�4��<�W��{� �ak��R�|�
��q���)�o�P��N��qnU�߽�,Z��NSaw+7��s�)1U�K����L^ָw.�]��/7��޷�7���w���䢤��f��81� �}Ɋ��k�{�~���`�*f5��D�k��a�-�y�KŌ@x�T��o���^�G�o8�I/�ʒ��4?&� �����b�F����V�9��)�[ǁ�PS5��C_/���b�^�ߦ*1oP?Y��8��g�N��o�5�9��Z~`�-Ȃ񖷏d�ܰ��F	_Q�92t��L�7�����}���L�{9n������Fs�	�@-0�!���pN��G�$`��p���������WR���(K>�B&�79pj�#=˫�fؤj(�}Pg.�U��G�}�8��%�
�Fg�T��<D���Х�� �"wKvT&1����T����d���л��^W����~� �e]���ܙ\iǐ�<������-J��J��
�^�w*xQ��sARK30%ҝ�����FH+�x̌G�x��;09��G�RM�42� ��!����*3��Fp����D�f������Z�#�o�Y]6qI��(��o{�߆<�?��3~\�Ʈ��^��"Ք�G��ܽu{\($p�c�c����+�� ϵ�t٧N6\[��I�G?�-��v�t _3J�=�O�-�a(����BO֧���ú!����ѩr�`��Pf���q;G�,M�Cb�o�@m˞�C�?��VCi%��Rwh>��h�y\uN�����c{�,e�ZƗ���9���B�Y����t�$�J��O	
�azs?mY���/e���%*���=�c���������)f��tR����Y�7���0���o[+.s͞���U��=2��ƀ��Lǟ��x�:�x�)^,��mF���s!x�q2_)T��\�s9���iP͂&T^18g���2@q�E�Qa�?�Gf�YH��(z�yy�ݎ��m��Q��4T�Y6�\Y�����8Wb���wXp�M?X9T��d�bQ��BFL�']>��Z g8RB��zO�c���:��I�4��T�*��'}c�"i���!��tr�#kr�W^� �<�%��N� ��_���9���&\�j`JJ��^s,R��3e��6��+?�.t��jI��9lk�����r}�j����+^O'A{�
=[�ޞ���gj~2re��=��������5��w����ˁ�]���9npqm]F1��%��r���~����8�Ӊ2��4ם�<R�;�P���P�_���9�d !�j�.�T�3�\eZg̬԰��P4���[#���@\�B���x=���O�LA4E�@�B`YMX#��'�n�>�ds�wv{X97
h�?͛\rm9lxFĽDfo�����N狯���y��k�����*H�$�T-1��[R�	��
q���>������s:��W��ș�_��c�DT�� 
��'�@k���:������?↑x�1*^ �L2��;����v�7(���ތ�:�]��[�!.��m��[�
.�)�<�F�!���>i�X鄛9� �V�W�j�ز�2�?�˿��)��DG�b�頎�e�ɤ��!@����0qi���O�rcA
]�~� �Y�s0���аh ���QAUʞ�$�9�vi�Oy��<dj�c$u�|��*q�J��^8���º|]�㪇�vq;
S[�Fp�I�$�7j���yX�_{�h���/�ϒm����-B� B[ofo���KÎ\L�9%c,{?���"� X�t$�Lȣ=�J����ݖ�c���$B��9�����3�7Z���5Z�MfF\|1_���)`7i-�h6��x+Y6}BŶ���t�^�/u6>��8�I1R,�c �r^��qIM��C�I�v��`� �g���I$e�IC��ɠ-�~�LX(��WS��4��!W�;�����#$�
	�W&�'�c�!0i�J�}&��>FKI�JйuW^�{���*v�W��H��X�x���FHC�Wɠ!Q��a\pO��g�T��P/*�\|����8������ ��ץY�g��햅D:���2]�!;��t:Jq�>tѫ�&d��L���͎5�\Tl	#K^Ƣ��P�_�xK��C;��L���[�N����#����i
SA~������Y�[�S&�V�m��&�m�܋@r�}\0�Esi�4�@ă�i��X
�Z�VFI� kgV��l��G�z�'7�O���Xo ,ׂ�S��q
'���`}�.i���<��dTã�����y�RjD��Qa��z�k���:���y�T�(�����^��zz���4�y״�!�?���vq�@9E
4�CX����$�0&O5������4&���]���"�݊�Z/i���B�h��9$O♀ �N�u��V��A������(U$K�$�d���:��vY�jQ�D��� .k��E��ܝ�� i���q���L�z��~N����� ����ư���r�yE	
���n���[r��v�!�	~ �е'柮\�n��]M���#n*�
�t�H��V�����l�f�g���2�ס�ʏ;�znH�;~���(���K��C#�4��,W����� U0F�4���:G� �0I���/�t�U���Y�����DM"��2Oc^��,����p�R��9[�}����Q%� �Gv�̀X�6 /�ȅ���
BU^����_<�Q��5�+%�&�Cw��
�16��2II��os�
	@��ꊰ`�q��K
;3�(�d���5�2�ay��+����DNC���,/E'���K(Բ:�.,���#fH>�e�Ϋ��Mr���'�_�1��m��}�~{2L���u����ېA�����p�妺�d+[���jP� �6a�e\������+b���5��܂L�W���h���\ �ź��-H�J7�����N��R��>�43:�z7�s%��pN+\�ϫ�MD�Ca}H�q�S�����#���rV+���b9K�;��2/
u�Nns��R�F�`Ǆ^���O^]Ī]o��zV�/�I�ӑ��ᥠ���"UOQ[^p��k:^7�2F�__�RE��ۯ-��[�*�c�[kѴ�cB�Z/ȧ2�e��v�BÔ�"������"�>L U���;�Fv�(��O������!���k�Z�݊.L��Y<�j�(�Y-q��'�b䄨�6��y�R׺ ��q��ĸ���$l�,��9 >����29=��;b>I߯m�������fy�!�r=�`�9�$�kt�W,|>�P��/��[
x�P�r�����&/K[W� �1�9�h(�O+}����N饃7��#+���Bw)�%�gQ%�H��#n@ޞQw��`���5�e���ƥ�ot<��]M6A�"]Yg�����͸������P[��*��x�؅,(��'��밈X���:e��0}
5Ukk3n�Cop����Q�A�uɁl���ݚkv�n�D��h^�NiT�q'X�J!Lf��i�<0�
��H~�V)�;j&�x����ŢLv��~�Kray�~�ٷ"�#�ڶ��Te-6�]�_��|uAa��w��n�\L�?!�	��Ůzլ��\���Bˮo��#Ё���}��N|x�����wɈ�S)�i X�~���>���v�8�y���.��H��"��~s�.�FK�}`�tT�������@h�V������<�{u#w"p����*Q��&���~{�����̻X�s;���F�ndA��g3��F��T�Ҧ��r�~�+��]:\wo}v���8B�[���\F#G�P΍�)�q�n�\�yݬ!*H�u�w�h\gvd� �e���L
�ĳ ˮ\�5Y���Y�����>�v���/�!�r׊�^�
��C�ɪ�Idũڦ>E���,'���Մ}��ֱ��t���Q�5�Aʹ@?M,{�^p����#2t�Ͻ�Q���ʇ���4�S�$N�j��}5�Ɓ+�Q��P�e	CDq�t/긴�>>��P�}��sXy#�f _t�R��8B�l'E��� ��xN7={�zmY������%��;�`AC�)�H�Yq�I�l��(-�OFqM�� 7h� �b��l�x:/^�<��D
U˄�|}��	��Obhku�-�'Q���N#�r��( ��/ֹ^Hג���X}h��G�o'K5����PC�3�(~��F�v�k�o��t��Ŝ��Ѭ̓6>���{qM�d���MF��y�V�K
�4���:��&�3�`�_�����ך�������}Q�XSTN���ڗt��cf�|��!����f��#q=�
��Ă����@@��&�Kf��?ŕ���U�8�����M���jU½��m�� ���y��@ηq�z��w$>�t�f�i��T� &��nL�_?�d8�\�j ��%��I�T�Nb��u?iI���2]��ܡ�{� ��BS9�[����W��K�;O$0�����ʥ��b���r%a���~ל�ݾ�`$a��Y�調hܩ�ݑ�S]Yǹ#���y_�IG;�J����EkU������
Wj6�yJ	�׿�
s�{s� %���32�Z"�x��ն��	�"�Z���lN�w�"|������2<Jy0Q��!�ǯP�'6��8q�}�|�%�o߃o2�������U�Eb:D���k7��do;�{���Р�垳�y��K����%)xTD��tI��>W�}J&R�F;k8�}!}|�9�I�)������$	��Vb�W�gJ�f� ��.�tȫ��Çy��5)5�ތ��֊-E�[B�CJ�b�c<�M����hY%D�1�E�Q�ly٘nHs�6N�FLW礖ff~����TI�Ԭ�k#�#(��Wr�?N7��nz,�M���*�KP�5
��6*Ꜻ�b�J��`� �
���aZ��[MZ�H��հ�d�����C)DĞ
y>�xD��30�O�.�y�CȽ����b�lx��3F��bt���)K���>OjEN��`�ڳ�����A�fIΓތ��$�J�+���g��l�)W	.�����&������wVȆkT�/�!�[�7}���	��U�m�0*1�%�я��J��A�����ŋq�3r/ӳ�ċJ�{� ]9��c\$�j�^mzf��|��.�Cu_)XœY�4A]Ӊ�Y����ڷ�\AϴnWX��2������j����Im1k��k-N���'������[���� ��\�sk��hZ�Y���.W�BP�UQX� `{Oi�v��5�J�e��n���,�X�V��H��u�������\���+��%X!��з����X&���
Q3�HzF��9\�(4(��uT�DG���ɴ��:�G��"`��f�tL�sn@4�����8U��LT6Ģ�V˙Tc]�m�����7�4n8"pޕ��K����эT�q�%لÍB�"�9�#�r��H�P��޴����b�T���L�"v#~��1HŰ�2��^c����c�Os,q6��R �����e���p�
�v�n�J���s���SES�� H��Q�,\)�h(�j1߰<;7/�	�O����֮n\���c�����<����m?!���Mۤ#����W�3�Y�y
6>��3����?�u*�@r�v� ?����(أX�xG��Fw�%�d�����`�MP@m��v�pr���[���W�B�h:uۘ�Rn&-�u��Ǣ����Z��+g����R�*�ĳ��9���W@�w��`��D�QV����h&K 1k3���*s����xܓ�5fGK36?���}ֱw�-w�XDm��GU5�M����W2���l�I���991rZg�����iL�tV��{GY?��ٚ�N�PU`��sq��mB���%��)�T��:��>�f��N|�82P��>�:��/Z�a�x�	{�]yU%T�{�틺�ȑ��p�R$��]��V�@)7��Еk����_GK�:�S{eDmB�qAx��lae+����XT����'�n����'����Y"��~�'��s�� ��4�Ԑ?����J��.[٢�hc!ŖGG�:>���\(�7m{'�8��ҫ�K�:��K2��r�Q.J:�j��F'�AX{�i�s���SnP4I��桀®��*[�G<!���}T[!T۫��X�����2E�&�N&�p���߯�iR�Ӝ%T��
F��/��Wͣ�il�]����EiU����q:���TSv������d���߽�>4�x#U���x�1�vC�i���%l*%�d�;���,�bOh�H"Um�?��K�3���(���OS��W���_�3��7'!�Q�6�2�}wr�Ն@|}2�U�L��&�����^�܉���o��Aj7"�e�.,KϬ��L
c����q���VS
q)�\�R/��m��Q<�ݾ�Lb�&>�K�4ݩś����E�{�`D*S���T��3�T�π��̋� |�5L���$�B�U��~0Rw>Gqơm�:�ժ����7�E��h'Mӷ������`�=q(�m/$����ɮ�lu*H��b
Yޒ�
�.�;}}��v8ź~n�/�LS.�$	��D3��eֿr�h3o����H�m��D�j ��vv�I���ٱ� .���4C�4b��g�	ǒ���\3���ڀ�!��B�@�=t�Zn�����K� Q�І:�	�����X"�	"jn�m����4�-���u���M'0��jG!�0�0���MC��[�뼿��X�..Kl�����"���=^��|z��B��}h
�/V"s�P��>�q��)0�]�ZC��2�|0j��T�g�І
6Cp�DC��=[f��j�Q�S���:��a>-�G�-;y\<_��
��|������W¡�7ı#n0��kSU��	��M1i����+�d��)j�J�� ��OXy��u�x����?8|u����Pє)�!���s�濍��"�L�>y���Y:���K�DD[�6���r�m{���>�z*�@����
Y5&�o��E���� ^�(B�m��[YԼU1�	��Q
�����'��d{����L篾켸�(S�CB�En�V�|p|�c0A����8�E�jBEV�gsWa�Ӈ������ǹGx�(}O��O�~�(m��+V&N�[�����O�aY��4��M�Y\��ͫٵ+`���o�l�;,��>�!5�mK7�Գ:����[���)3�![��i��:PN85��_�J2��!xj|�D<�Ey[-).�?K$��xN�p3fK/�(���uw[w���f䒆�l?J�}tM.��:CqI�����+�|R���_��,�{܊l͚�e��Ղ]n��പCP}"�ߛ��a��b��4��~����1w�����ˈ�^�	w5�p���Ae�t>�/�c9/}�\�c������4Z�b|g�'�	�����Ny��m�+c��|).u(�K����f��0/�����5��<�]���A�q^��=�w�}�r��8�2��x�mV�wAيi!
��XBk9��v�������moF/
b{WQ��_��C�Ȅg��"��> �i;�dEN̶<s�j�X��,��hSL4�}��ܿ����N\[
Ck4��˷*���B �a��ynV"wK��Ж���$�Aa�iy�Ӽ��
&�d��UIf-���w���F�����!F��=?}3�6�p� !����� ���T��@��ȗ��Ì{bl��ۂ��4�y#�r�ܓ�۪�/!�;��i�[^
|V�;�X�Fn��/��)P!>u[�6/t�=�p���Z�,-���Bs�x�Cc�s7�>4�lpN5�����"&���
F48`n�pǚ��&<�Y#6�K����1(H�x�5�`H�ݎ�g��,�+X��G����VH�D0>fp4�%�AWzy�n��������r�`��YH��l G�+���b亲^l[Ee���~(�
�� �6�sװ�Mݮ���	�W�cJ��ͦn�b��UM��)�^L{)Q�~�(*�¹>JiX ��<b'(w�w>�x�i�̸�n"����6�)_��zX���(�=.<�����!݈њ���ղ=��:V��BA8 �3>��>�q�$�|jS:٠�z����I�7�1|��{��l��D����q@ӷD���9��[ PJܡ��p���g��V]��!�0Dp-M�5������U���<c�7�Ji;`<��4lt��A�1�?��Ȭ}�h�����ttY��(��BD
�Κ�H�\�����Ss�� m�i�}�&׌*�h�3l[P�dx��?��{�6㩟�am&�ǖ�3���ֿ��r�)�׶n��4�n�a-�q�n1:.�~օ�6��crg�$(�L~��O�V�g�%��PFN�ٞ�$��OH1�ނj(*�_�S�F0���l�]�u$�@(�Bu��gzm: ���U�V�"��.s��h�29R9l�7/-���c�F���	s]xb��wQ���e_}�����AG҃_I+�����p+c�<�ɩ�O���0��QLTܘ�k*���HžPv)���>�ѓ����s.0I��!+[�ҽO+��w�x[�8D.�Iy|[�˰��/���[����&��:?����q	�7W�&��Z��R<��f�ڲO����c�{��	D�)�� }u�2y}���\T��H�*z1z���7E��ޠ���h���w2H�)L~4�����:*2���*��0}����.[�$e��y����wK��T�^!1��>o�W���ٗ����������(3�IE`}���Ť��5J���NXA� �Gh�w/�y ��r޴:��I\��ݎ�c;��T��'���<4;���]{I����.�sb_���=����i�(��M��t�F��W|�TjOEZ�4d�/�7vm�jZ66O���+���5���p�p`0U�ҌiH����e L�݉d8�	��cv_��UL��D\����\`�(���䳀lwZ	��u�9o�aN�i�@�p�7G�-���w���[+��#�w�&����h��1�e���J:�}�M���Ք#G��+G	]}(yd/���}�П�#;t�W}�A�+������b�s$\��O�Rf�*�*�O7��`�	��q�B2�%k� ��زo.�b�0��v�X�������B�� �4QEp!O�>b����-���nh�xV�.�!�T�qT&�.)M)�����u��Y��z��o�,t�����-x�O�(|&x ��_p3��x������#���yO8�Ƃ�%'��`�������r
����lz� ��Q�˭ϲp��/YᑒW_�H�
�:;|�ź?n@#��6/���Qk&jI0`���k��&��ƪ'�u�n=�e���!7w(@��E ����BXh�Gl������0����9CKl�XEX}�hC����������ܚe)J���?қ���H�Z��<$[�X[HËR���Ęe��Qd�r��{n�r���Q竭��������*��f�
nm�P���o�$�¬fG<��=�6)��%2+����ApU^��+\d��Th���LNɭ �	ɦn��=v3^��}T��P�a�E2�3[������]�"/��1y-�QZg����UV�]�p�r�1��|#�L�T������{Cu��]eJ�i�8Õv�ǋ�v�n/��4K��H�_�ې�)��ǯg�Y�{M�w�E���g�X;����ib�%w�MA���ak�An���dvMջ�=
�z���AW��L�'�I��o�������ԩ��h��C��X�=����68m7��/x�[�[�ު�7�����ܤIU�ʴ�*�l��s��v��i�OL�*2��	%�q����4S�T�e��:؎ֳvmQ`�̳����F�7����fVa<���׸��ޚ�?��H򯿱l���d�S�V�j;�5s.�9x���VH��[�չ0���[��0_�m`9��$�[��T�1��b)��xH�� �
���kv���9U�$��ºTJ�1Ljks)AV�:��\v�����.��.jG���p�h/�]h,�0&w*���i8�䖈���ϝz��R�"<�~?�5����"��j�iҶ~��|��
ю��ᇻ����ݵ%乭U4�#�H��A��q��4�%3?h�4C2������t�,���+#���:SO��U�\h��W?�|�% ��3���a^oP��y�f����`{�4�'hƦ���'g�-:&��'��^���O!���*�G�C!��� �+<�r��o]�F�2��*�|N}}��Q[�fv7��"s��H�r|��NS4�}�:%�aP1Ц_'�P�������0!��;2�uR�f����aib����kM �$�)�0&h�S� 7�r$ˡ��$\%�#�����\�k���UW�#W(�O`�;o�Qz�B��`�W���%=�3V������L}K��$n�WN���Z��K���B�g�D/�X�2��>�2�L)�5W���M�d���䳪!h��&R8��O��m�<RqߕL�����G��&Z��'��9i�3�XV��mƱ�[J��KF/���E��78��\h� <H��K�˕I��H��2z#ǈ��V�le=1���D��Ń�4)7v*���a�k�5�X8���uq���[��.�]G��:����1�܁�07	��lP��<yQ����2!9fsYBk����j����{S��4{�`֑�ޝ��[u�;����'���:@?z"���,K.�����f��~`=�+o�
p	�@I�+[_��ٲ�� N)��2jxh`��{'#�e�e���|E�`!pU0�k.��oH$.B�뾺b��+����`.p����!?q�p�T���[��u�z* ����ͮ�g���>{�]�h/���NU  ��S�5��S>~�C�D��-I@.��қ�L��t0��0�*ɐ���s�a����X�,Σ�[_��m�����돒�h�Y0m�����mX�a(OH�&.�+�OpҥMZ�_��	��y����	��ϥS�l��p�x���0n ��i`VH�T�պ�}$�.d�xf��4�]8����u�Ե�Wt!27/��5ؿ䣊�@1<z��ÃS���R/FY��X��K�j�B��QI Y���C�W�>�������(�Ŵ<�Z�D��Wk�uDD.��}%YRdn&��/;��B�耭& ����F3 �S���$�[� �#^���L�}�������@>y�c�e��q�d�.@�Y�d��V�\1�@�v4�Y#��1�7(܌���-�ݏ�L��<�n ���`��e�{�"y��~�/T�:�����T<�B�c�7���S`��)}^��0f�Ԁ�dZ=����>��Y��t���
�lg�h+�`��~�H��$�|��d�~\�H�nIsyC����p�E#��P�>2v�[�׃�3	��T��k:�"�ީ�}E�|��1ބ��g���ɋdV���5:1q�;�����l^4�h�-����e�![���E�;0�(��T�03��c�0"��J��jT�n����^�O���<���6�zT~0�����*̥L�`�������6���w��b�,^��vt�J{� QQ��h�	�G��#��J����^�@�C�É_L^ɓ���?��(d����7<��)A� Y���ɫ�b���߂@��,R4�3p_OF��H��}V����Ab�O�5�tx�'cП����h\r� ���>b�	��@�w�@��Ty��f��:,�]��]�ّP7�ԀT�A�6SW�>/g����j�N�&Fl�
qW.U��FX�8���m�4|���B�p��������-��.!J�y*>Z�#n$�� ���hCH7A��i�Ϥ�� A�����(��wό�l:�c���+�Oǿ�%R�8ݽ�V*DLY��1Y#���u�/�zn�T����}�T�#�[���؆�x�s�����]�A|�I�y!GQ^(�S/��n1��5���`?88�[������P=�_Zy�c�`���*�ֈ��h�!�>���z�ߍ�Al�P�!rq�D�/o��R�M�`�0��bH�ɪ�#�y5d]�~�G�mLrL�:�3K�bk�0k������$��7���˟-������������Z�`��TSvh7s��br�
��k۝�)쟿^�3*���N�KL�
o$q��xe�=,u��zF����lon�@2t�t����65���Ҟ�]�[�5�(���{�_ W��u􁲙��"D?�]�w<�歴J�b��l�+j�����|u��1v@ѾN�����ޙN	����k���<���S�ϻ[�CrB���Rj_�zt}E�߫8��u0�*ZR5�E���^y��h
��+�l�DU���G�wS����N"�K���Jy�jJ���(y&!11vY�e�>	�a�s}Z�WF���g��&���Մ3��6"�^�(?�1ףl��<?�3�ӥz��|2c����ȣ�.�9!,�m����o���<�*D�������?_ J�u���S4�X�$xb\��W������o\�a������#�X��K���T����~�!���?�Du7o��N�k�u**�'�$}��$�'\�	9��8�Ǫ0J����ܭM�I,�&qc8JV�n6�ᮢ��K����]Pi�5;Q���$����S��������>��y<C�+]�t�.��I�>�C<��e�O������j&�ћ�\�#����a콃��l��ͪ�/�R3ܸ���8�0��D���F�vp%'J8 e���eErH��D���;N|�v��1/R�qO #X�==��ּMVៗ�2�dx��re�
fDؾ��^�:�0��~U����硣�oU�0i���4�ף���G�uq;$e�C3��C'�X0k���ox����]��	�&e)zu��5ZU��V�����6Mx`|g5ݼ;���:8o�Z�簉r�o5Æ����ROg��"?U(���^*t)N�TȬnT�K���'�\ō�y{s��������x��p�~I����Nϑ$�S�}&�'�"���?�)����v�؟�f%��W!��L�'V5����C裁�0� G�[��:�G+�H��(` �M�Ԇ�/��u����eF�$e�/�#,W�x�IqI�����}v)�PH	�]��=6�ua>�$��`2��A>I��"]aɡ�w�����PE�Jʟ˾�s/
� =C��S�Ac����6���2~6P�:d;��\�z���$��X���as���;!��I¬���s�%��x�k�&w�J�f�	�9���	�Cm��d���C!�$��r���U�`�v.H7�!l �^[��%]n_��T��$�N!�&Ģ ��*�:j���'���6B~wAB�s�T]L5�*Q|�۱��)���D4?�$bH�߻�G*4���{���(�6��y��Ц�\A���?|��/)��>���@��=\�m�L(Q>4t{�$B�O�tm��@�&-ɐZs;����C����I�$��N���t{m�����@'��E=�T��8�|�~�Ԕ���/�e��TZ/�U�0+�����,e6	S5�$r���R	U��#>F��?D읡ОN���ct*_%⭢���0�LY�VaŲ�t�ɜN���a����gŎU�I���\(�E(o!s��3~d�v��^ʹ���sKB��M�(��-W���G7�w�b=�����rd}Q2�5hx�{��P�3�/��^37X��8��eӘ�X8�D>����\�F�<T�R�)S��W��6ZG���V�N�2���f��0Jf�ӓ�d�f[j��x:}�e"x9��o�-�m��H <?( ��l��窾��M�~��ℓ<��hʅi	:ߋ[�MH��y@w��j�D�	�����܄���+��2����)V5�c�6�1h�ߺ<+8��d��/��U�>�C��	dݒ���2��i���v\��{�E2���hAkg3n$ha9��u@\��i�`���C�{�~��:/v�p!��V|95�Zu�R��*����fB�ʈn�NhblXEߏ5r�>�0�N����yuЦ�[5�ĦU��s	�jzȁ��QȔ@	�leAk���Ք���E����C�j���,+X����ѺC�[Tؘ�iKdB�F�J�s�|͐j�AԴ�A�/x
Ѿ�΢��Խ2������'o�+_g����r>rf���K���G���`��'ud��rُ8 �֕��=`�?f�
CH
EA7o��m8βy2�u��bt�j3Tu�2*Fo�mc*�N���`Q�NᤡBfmk	�ZmDunՂ��0�)m��M7կ�	������k��,�S��(��w�4���W��0���. �	r3jʹ��x�#�D
���݆�:�V'�N���1]9m���rd���d/X��Z���I�m}�n�(�PF.u�m��/b��.�o���+�-u�:;D.p����'O��mB	�<mk�E�X��N-�%��~�_�=y��:�D����[^�_���)9ye��w�Q�1�Q�;� vf�,�b�T���o{�?[G�L)s��kp2�6aϓjkopz��l�֌y%����n%�T^Т0h2��R�S0�S��I,0y ��M�ё:tB<3�@3�bv,[�l�4O�	�0���c2�G�W'SÑ��"�1��#<s�"�����WBF}���m�yp}�}Y����!�_-�+>spBya�+�G�L����5|7��v/-�#�́��q�?��!\� F���G��胻��X��~�/�^�ܱ��n��CP�W�]Ãe��?u�u��a��ޫ��i?d4S+o"��+�}��N��d:���Z��@U�K*���NQ�b��勖V��R'���@�U~ �S�ުN{}:P�B��u�C��gN�!I
���w^��uV��)�	�q����t�M�"���t�ʽH���ɗK�Ny6Ŝ1�k�'y�{�c��P����U|��ɂ���wGࡄ)�����H����h^�~-gk��Y4��ʨ;����Q5�.�sΊ'*-�F�[��t[T���=M��Ң�
��C��{s�L!Db� �i���9s�̈SH4�_H���A�e&uc���]��]���W��x�:�I�i�"������soN�T�M|/�۔l���HX�_�����,I|�yQ:�5��<H�X�@�D��B���nD^�6����򫊄�ڣ�m!��[������[��%'�^�^�U�]�S1�119���-�IXj1eGY�P�K~�p��^^���y��d����#��@<��<2�l�y��;,Y_��iq�%?qiN�o_\a7)�t�k�������+�P{�ђH4���5���J��H�I8��P5�����	_��)���"��UZĻp�J��z~���Z�g������|Ň M-A���^R0#+}NL���'�����}��@3k2�M|���C��ۮ���գJ�A�vh�nfk ��
�ͳ�/���Z6ֿ?�e[=�_��:���-Vʤ$]�6����0���PT=�KV�+�d��;��e2Ql�t���	�w����y�-��;ns�x(�w1��B��Կ�mص�a���i7��X�Եz�.̬��G^�&EF��Y�2�����;$�'�q���v����	g�=��Kq?��F~����uqr��!��B��$���"�_�<�q�P_��S��dv�� ��2}�0�a��fO�VZ�1�|k��4�B;�;����ˇf,�cK���a���ǹebk#M�g0x�ϖ��C�ɿ�;&PV��d�����p�~`8�e�'�����j��y�m�ϣ���)��O��� �H�ѿ桠�v�,\`�����݉U���1�,9�H��A��m7N7R�����)�	V�,lŋt���*�?�y~/��G����/��T7�q�tU2�bG�z���V�+f�ދ�@�V�*���
{�Am�ֶ��5��Pn��G�5=^� ��(���%���`E@�z�-�
����˜O�������Oo����p�ND�2~�Yu?B�l�����DYH��C�Y|�w���m�r2$��e��R� I���Cv��-��ԡ��jZ�[�2';)�����	����TIUr��Ep8F'jDK_j���H�Ez[/C��>�K���n���Pw�&৴�8���q�ƈ�%�	]�#���$.�띩��v�OT�_OO�L^{x+�hR���̡4�/g���W��f:���^�b|i5�B��J�@NP6��A�^�Fb[:8�P��܈����7��@!7�"�}N�#BL���}3��:xݩ�A��zq�'&�>��@VS\�Ď�{����k�;_�������J��P��'e~��b��5�	�}���z�P�W��AQ�؟��@�&����'a��:�XZ!�Iy�{͊��>hd���+��W8^;�!76�!����Y���]?#�Z�'{�8�ܥ�gV�w�����,Ki= 7�.�uR�F�Y8�4-W��{*/��;Y�)�ɸF~���$�����9mR�;$3�s��+bO���C�-%�H�m]!<��G#���}G�k�҃���@��S���<��\y,���o�+�/Oa�Z�[�*���vjw9[��c�I��z�ө�/�82G�{����yp�f-�	{#�6X#�1ӷ�6=�T�K�x�����X�v9C%5in �B/<7���%К,��Db��<��]�)�6��7��V2b/6���`���f�оY�i�������=��ߜ�%��T�2���;9�Q�l���x��Y�$zb�~���I��/��Jh:���'����>��蕵�A���<�8�fx�K_���P�o�)�JrE`"�An�K�t(��9:���xpp6V��,�91B��	�B4�v��.-~�}S�two����ʢ�����uv]ߣu4Lz46{m��}m�f��`�~L�e� ����ZO�̤$��8�>�F~?�$�h%�N��[Qt�8�h�o?�`x��%?�z�8�P	�HF��7���:����$t������&�6���=0~6�#e�1���ѡO�2�:S����OT��_��-��?��d���uwD�3\�b����Iဦ�΄���SpnY��H�%��;�l}^�t��V����P�*w���]A��I��R��H�>!_*�`�1.���ؐ��y��J������w�Yv�ù��r�6B�X���dB��n��	��Jv[Yp.g5� b_�a�J@��q1��3�	[�p�EiF,���Уѽ/�`������]Eʬ�,#�݇�9m�օ~��&Dryx���hyA����_@w�g�fJ�c��k�/�Mj��8���R��������c��������5"���!*(f��\ՠ��y���o|�?O�i�}ߊ([
%�A�X�*�N/MǕ-{^�4p��(��(�� ,�d���lf��RuI��r�"s1��1X�c�&�������1$��x� ��&"͌b�?=�����q�5?��9�z@Ō�nvc�#�|���D�߁2L�R��`?ft�
����8o�5.br����Ô�7]0��@^V�mMg��8�NQe`
3N��a�N�xxd��Q�lC"y��!�@7��Slr�;�e�˗̓A$��7X�xlf6�����&����A�쌤0��v,�`V]k�N�דǣ��"�a&��^R�����:�~x�_XaE�2+|6J�KL�	���#q�j�_�3hA���Q�1+]�T`^�p�ى�P˦�ѡ干�P�4c7P��Um�/���p��}���=W`5�~j�l�PBB��y� �Vpi�����ԭ\��}4�L2u��9 �F�a�z�b�e�9�|�xA�N~��.�`W�h�_�G�b�&N{X~�]��A�?M_���	�+�?����/Y\J*Y�zj�Ms!
�7�h_���(L�C"��,,Dm��E�}V<5�ԐMp� �E���u�wqc�d��rl��u�ɿ�){H;��~{c��Y�-�R�V6�9�^�͐��C�d��d[���* D�� Oz���z�*���`5�����n�8��_kkt�6V"�����u�g��mܧ���O߳ZTc�oUv�:�s�ؕ��Ͱz{P29��T`:�͕��.��#<���i��p�fEu�.<s��'��D�Q����gٜ������)��B�;��9kG�:��ɜ Rf�]@�-1�����͙p�Uy�
#
r��x?�~T����6y�ɴ �QW�օZ5�Bm���n���:߅����	�f���W��Q�|%f!x�_�}�QهR3 C�=jv`i��a�=b�MM��c�A���"�����N��\@o/=~�{,�<�%�l4'�������?k�V����l"+P$T�=�ɡa��2�пQ��є�@+&"�Wgu�ɣ����v9�O���:�A��0�d�Ɨe4k�u�
 �U�Z 0�!���~*�8nď���OE�VOԜ��4�4�.:��|𓠹'%x��mtk'�'��{l4�����#p����9n?v?r������ |P�1�!���A*�Nڀ�e r�$MW�v[�M�Glq�0x,L#M�����le�@�93�8NT�ؤ'�3$�����@z��Q���"�Z 	�J���]|)���ȏ_7�Z짫�t��G��,��ݧ���\�Sj��l�O��.��Z��Z��%X?6�:)�n��gI��S��ѯ�V��Hn����_�\M�L��I���� R��4'�ꉨjW�r|:]�i�ʈ6�D5����j�
��L����E�6Q��UZ�ӻ�YK��s��;�̔���*���_P�!�z1"��<��������`. Ki�>�<�Q�ԃ���}��c�6��
r&�ݬCa����n�Sh����QA�u�qN����������S���2����,���4vg��^�}�U�sB턊�+��RYh[[4%[L"��W.ܲh�F�������u֎�?�j�bެ��C�DW���\���Q6d�V��Q����'d\����C���$���֋�˃�b�5K��v��)��q �7�^K���c�������B�r
�
��y
핃��|�E󡁦zC��MN�����~JEx�����d�+��"rT�e&��=��hsZ�Y<����O���~��GM(���Ғvޖ�߲�}�z��aYv"G�<�dO�;H���!��jӅ��W��|r�қ�l��U �WIv����s�p���h��]SzlMG��~�=����bz櫾m�/���@�P����ַ�'dW�\� �ѷ����$��$vm5o���֛����i˂�a'n�uPN�P���-'r@���NDa�����+nKe- Xk1�sL{iی��5i�k�Y�3�����]Ri0���x�D��4�'���#��0�!���f�:��UT��1R�������֮Ų����ï���SXM٤,N��U��:b���D�7��bx�q�[y��a�?-��/3Z4�M-�q7�o=�8y��:K���%%���T�,�O�!�-0���7=��A�׎�_���B�ޓ
�u��㐧[@k��^�
�)���ͭ�S���0=�{KU�E�C�r��պz8����vEu�(x]�Ю�`������D���$"0 Ac_9��<���#���1��.'�dx�����G��6P=��!&�U=�N�U� [!�(l)`ج)�`qrs�vQ�5&��q�)31��E�� ��V^26e�vޔXw��KDߥ�Y�6?�.LZ���3m���k��uR[W��
��T��lOQ= ���ü̴JU^������
�P��Ssw!c}VGڃ�'�µ�'�AX�G�4��T�{EIu�(J��A�t�"Mz���L:�rXץ&M{�vH�7g��
:Ȫ�ի��?E�����eb�_�	��돛�t.��&��P�9�����(��n�����?�����A˄�0�i�u�t���p���EE�Ңfc0�W�1fM����S����$A)�F�Ab������!�r�昿`���[֘�E�Ϭ�R��gJ�`���p]�'+�ڽ8�(Fi�u?�ˡ+u�_�I�e ;�����	�6�	��QK'�5L�w{�;�J1�2��~�9'��Q��*��-����I�ma�S��r�45� ���$ɖ�?9��������>�I��Y� 7�o��,����⢻	c�š}��m�i�c���K��1Mc�uAr̨Y
%��~��������K C���'cY!S�>��ƔX�l�M�|�^IM.����˓�l,>maX�����g�9V��Z��w����5_eĨ����p���v��!�e��ϷF�검lBU��$�� ��p+����2����8�x
yֳ�,?* Q]�zhsن�a1��amͥ�f_e�<E�z'3^����/���s�n��%1���j�٫�x��n�I���P8�}��l��:�}'>���<�4ߴ���D�	e�$���\�Y:�l#���e���!����AA�$$F]��tq�	��G��(�|g��4����fN��Y�+��ؔK��Q�*Iogh�<����C��E�p}~�͵��&KDt	s %0u8�O�O�����Sș.}6j��͎s��}���&��\)2��v������|9�Gvټ�N���F�F�GyZl� Gٻ���z�ǣ�2�?�ͮGxz�P�m"fm7|^���Ǫ�xتe�Hݞ�
uXuJ����UWeJB� m��Ɇ�M�����Xߖ�f�{*��#VCj�Zu�-���9(��u"W�Ւ�b�2�
��`d�r4_��pW�14�q[�ӼO�md��/���Z�1u^������z��_���{ի1���	��4�2���>�N%���W�����X�Y^��Y�Èa�j U�0���2FO�X�&uO��Y7�&��k!���������V�cw,�G��,�D�'��Ê%8��l�e>F��n��:`K�J��}y�~��� ��%����O����-E��J	�t��J�贈/������2���nt�lc�tR���k�M�k��g�|���c��Y�	�{��*�DÌ�z!�R��>2�O�l')��%\A�_Ї�����@&rS)����7a���(���yW 6��v5rSql!"
d^�����X�O.6�&T�{�b2��&�*n39�-������	>'�ī�`v?��w,���P�Rw���">�$?\��C`����O�#�w�����>'�蚾^������z��v�(!���Ɉ/�Q��6��i�])��4ġ��FW��h�}6x�k�ϔb)��}޹Q4�n;&��@_��,���Y"f�dv�s
x.1t���OR��b�f�i�V
Q��ͺ���d��9��R�`V*;uj��M�WRK��v�� ��� f����Q�����WQ�砩bX�2�i�;fd"�'�3����Ⳍ%��`t]s�B�EMW���B2^3��_��:��ڜ�����L�U�8}]h�ɴJ�˥a2��Oۋ1���p���g#Pah�7N�4:܋e:�Q����qu6����|��RC結5�zu� ;����Up�M�^���]�n���-�wW�j3~>Hjp2�����pq�2O�D�c<��z���z;�4b��@��_��q���E��8��\�?˅�J�n�b�:C冫�q�t�!��%�G��j�LΪt�9Ѝ}� |�ztCP!�TD���!��d�엇������	��wi�Ux���_f���d+�pP!5t���@���u�&u����B�ԠOB����Ԕ��T�[NƉE~��]��[f�M,d����2ү�e�.��~F��"B:)��Ԙ��V��v2،�BH�B��-�1w=�L|I)Ő�u?L_�Z1��2PO����Z �=q(�I|T��,>�@Q���C;���Kz����҃��F4�B��Y����M��޽/5��Y��U�͇{�/.��]�"�S#���-s\�ѻ7�0�l�a;Uv݊�BF_V���.�-��,���'J��9쾾�I��~j�D�LgTIs��@�m$���°ۥ��m\���(�ܚy��\�H~�~ě�]T���(���\���3P�9;~�"�4���5a�o�������
a*�h���A-	ځp ��h����$��U8��F�<��K�W����9���H�ε�k��e�����[�&H�˩Tmn�~#4/����:��Q#.��))�Xj��s�r'�O��S�rpE����-V��+�|zc�u�bs$�<�Ӱ��b�����6�!hΫ�|�	ױ˞�XO���h�x�"Bςf��~����w@cV�y���*�gBр�k��!Vdr��뽚�w�x{zj������kU$l����Xm�g1~�˨~B�>��貿�=��p�����/�J�BOf+���x�Өa�@)�&���+���X���L�n��%ĩ�wvf�pӝ�দ�d&a��Cs�	ѽ#�W9FFn��mA�$��/�@]8�5������}��v:��.��O�͉K��f�PG}l�{[��a���ӫ�j^��H�o�a�4�4�[c��d�׈JO*�H�z�����R��s`�Y[�\J�=���3ٝ��L��]���J�J<?��IQ��n�]P��\���	��l�����6[���b���_
ϳ		#k�&�߀#b�N4�KJe]N�� ~���N�p�<���+t���p�eOa�����e�Zo23������05�+Ly>��[ˬ�Eӕ�D��~�'�0t�)��M��G2�2��Xc�\~�0 ��Xo�s��&��]�t��1PV��Y݌ �)�Q��x��.8�F��h��L~�PqhX�,<ֺ���r�1�jW�{:y但��������|��u��A��e�L_Xa�׿A񱒢Fe����DԻi'8j�s�;�ʺ=�GD�����j&5%��� ����|`�T &,t�8n��z3;�AU`��"�\��o��,h�#�����ШÊ�Օj��Ӫ�O}Dj��*�����ԅ�CW��o� �ߪ�nX�6)� U �,\�ATg�Q)��y�-T�:|E�ؓc������6� =O6��f�^�I��|ȸ@/)~�%7[�o�1h�i�K&��z��L�[�pv|�p���+��{���
���B2�lH�E��]�Y� :ڢW��1�u�̷S������<گ*���U����Z��4~,R.U�A짧��e�xr��h���p�)����%i���h�qQ�!����;N�}X�h�?q)z�$o2N��?��l��ZS�E���h��$}WM P�sܯ�]B������5Q]"�x��A��jPpw�#�]��u?<��0�%P�����DUAA�G�H6Ym�/��ɬ����l/�vg�<pQ�=^��a��6���	g�1*���i��U�-/dJ��.��b�����j|��lY�5�M+&a<�C\|~�m����<�OY��<������;�G,>eK=:]u��q��o��"�~�� d0V�K�JQ9��f�h�!�h+A�
ji`��p�