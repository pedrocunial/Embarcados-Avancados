��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��l�����f�J�éy7�=7?�w�e���˦��X��(|�EN��:D�*��{-� {���hEې�_�p�P�Fॹ(����ұq���[�A�

��я��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c��Z#��5/m�c ���i男��,�9;"+_V���Mu>�*|���ғ�v�]��O�[U.�����Afݕ�(Ѽ�@ZL��d��G���J9刖�iR���-��:Z�_8<"Xg+-��ZfNL��m趡�>)ϫ�#;�e��8�,n���(k�~�e�ij��������O�նz��7/cD�3���&Lť��	2�� \���> �X�s�L�7k|��z(����?����dX*����������@�W���+��J��7j�#Hm;{�0Pzڒd��*�U����>H+Tv�f�k�!�c94�:�O���A:ոF�|��m��&�28�Zۼ8�@т	�=t϶�����S�PĹe��NVb4��jOЂ[sI���yvF[4C7P=��4��2:�+�$wX���]����+����$q�$H)����KZ�&�`v��:���蕅�I�2ݱW�D�/I�q����$��+Xk��ڴͼ� �Auߪ�4F��Qe�֗V���F)�@a�F�p��b��P�K-�w8��?���CɌnr*��� ��?ѓ���I����8��e~�f᥊����Vڛ�����2�"�2�r<ͽ�9��X�h���s�_���W���Z�9J�M�UW�Y�n �,�4ˌ	���hS��lB�E2ꬻ筕���L&>Լt���J����$� t]�b��'D
E�4'W��4L$�� c
��w������r�\�ZN���+��p��y��FuU��2���gq�T��?�xImS�U�@��g��0Nܑm�� �a8>F�mIBRG�p:�T�yVtu �Cn`>}�d�2�� tML/_١i�?�a�<�w�*?Wdy]^��2e�)��0��;�	K�J�ӽ (3! ?/خJ��6'�-��9+� [X�'�{2�f
tV���MD��Ղ��Ju �, FK̫��Y�셽��
�Ơp� ���-;�l�譀l�L�t�|����ȶ|�p���0ݓ!U�S�y�U���0����H���X���|�F���V˲B����(��������'K�'�ǅ~g�H!�*�&����	?��e$h��w��o8�}��w�%WR��Ak$g#e.�6�^�vh�p�G��C���7���a�}[|15k�L`V&;^ti��D`���&0(�:�ǎ��4ڥZ������؆S�S��`���I=^.�4�|�[7_�<�����F����&���RE-�S☝ɖ!�K|+1�Շ���[ f�)@E�����CQ�nC�k���T`���؛|	cM=e�2�s��!����|xY�H2�:W�Q�C����CJC_F��D���+w�"���F�
U&�٩�;^�o�E>M��لz�w��.�/����Q9P��Ǩ�|!�Ħ~[�]
 0��bP�M��>�ˣB��#hs�-J�ؑ�n�����7��n	K�� ���N6UG�G�����IӐ�+���<���� �V�}��g�R¨I�R��$W�*K9���,4t\P�@F�Z*lǿ����iD�@��ZFd�{?ʯ�!�)��%P�� � F�)�,�F
A�_��xu�<��I��"Hm�K�'$V �+�4%44�n�[�۫�A��5ʧfR��b���ef�'�?�~�b1���S�۰��M]SE�����k	&,��&T�b���T�>5F��^�/M����e�V��oV(Yh��Ь���R���P]lYt�Y��*�������+m-���=���0���@� �1��=��Ud2C��}�����dn�(H?�E�)�Z{X���(a��9�����a�d��jk6�n^g5�|_��oy�5Դ�^�}����"�Nt�H#�rR��EQ�@>�aX��Ҙc4{����U�B���#=�):j�:�k�";I(��%���#�Bg@���[Z�<u�,�4Hg9!�U}uR���b+ U�(�bH�x�����)��j�rT�� I4G��a��5W��3\ƍW�k;L��_�%��|���H�w�e�UL���o�>G��n��b �i����fY�����'��7��N(�B��@�&�iZ��"K��_��1�c���#h,ǛAd�R���5t$A�p��}����&r?�0�:"�f��ұ���h�*��A���th�Ԉk����A���}^╢xG�
oejb�b��S�ǻ5Iٹ�S�����I(����tc�H�N�I]���~��AXi�T�U�|���O�'\CP�n,���]Yߧ�ْ��WX"�V2��j�=�kTL)�A�sP��*mA�I�y%6��
ؗX��Rz����z"�w�����k���g����۔�2/@�$vl��p���ƀ�%��h�G= >t��P����i�B��V��Q�(�d��GI��X`�Q���<�[lU��&��_O!#Ah�������΄D_mz�d�K��Bt�j?����6�Ԡ��f(}t9�/�wXNd���jӢG-�[g˗�{9F��`�`S��Χ�E_�SJ�y)(íÎ4�*���h�n�+���+(۔զʏ����A"`r�����1��i�O.n`)��#�'d�O��� ~I�����̾�f�/�L�c�Ŭ4�7��9[�K#��ǹ�v]w����e9-X�ׂy�Ml��6փ���݊�5%{}P����J�l�KU��6��?%)��!.E&��0px��vUA�x�A2��Ka8#�F�L]�_<j�T�q�׎��ǯ��i���u���ǚ�J$,�Ȣ��,�
O���$lՍ!|Q�\�O��9���^�
����]�#x*�53�3�^�$i'`��X~:p�P(.[����
�A�������v�x�Y��	H�_����[������[ܡ�(S�a��`�66@*4�v�J1�|b Kl�&ُ#5bt1~r�������`��yTWp�2(n�����G�����o3�#4�~�����C�@� nja��M"(t$�߫�5��?����0�s���-N��k^�=�j��&^vzR��ʨ�mV<���P:ێ�7e�FP
R��gV�<�êw��l���d�hRG���o&�Eڮ���P) ��S>?߿�̐���h�WOjl���~�� �d�������e�sm#�t����v��_W�:���#����<Fu&�f�>�CL��/fP����W'�m�ڡ������-(���Ƅ�0F�]�l.�����F1�F��n����1	N{OJ��?k��G��Ro��5���X�h���	ME�[�[����A#�����9I4���̫Dȍ����U� �͋8�Ί���G�L�i{<�r=`��^���Z �E��
�WUSB����2J��[��e�m��8Ȅэo���*?z�,��W�cB���el�����1�R��2/�ҋۯ���V ��L���&��1���h����~��h�3;d��m�{a��_�����#�5�����DRw��c��qh��{��` ���z�᫮B��R��_\� ������u5c�9~e�e��+Ū���Pk<�v�s��"��͉��g0����b��n�B�j��.cg�J�E������V#��rQ��*�ߋ-\v]Z�c����Oe}&X �6���u���gto3����]3��P�ab��f֧���<`�*^���0+!'����m2�~�ܤA����Yl�!=Ȥa�7>���3��xm�@h,NL]`W>J�C�e���c�0s���� �8���]��41�����cF{����L�W��K��oa:.^4�^ytb�w(0���?L�C"��@9"�?"�^���Y�AH�=4�D�<�g`x�ﮐ|-���w�T�6@�v��(4�l�Y��)m�w�l�\5M�(�7�O�>6��Z���1���#�v&��$�)��q�v�V=�C���0�s����[-(�*�2�Zm+OyX]4c�GUzQ�r8@>y���9u���!җK�M6S���������M������w�w���G���$������ ��w��ξMI��%JHP�?wkU�uu���eޤ��>�t���2	�')�ny��+�c[r�ye�-�uD�]�qZl8,�S*)<���]�"�IEMm�J�/k��.7&�P�]���pq<K�T�]�����-#%*�a���#H���	_�V��9k��TD.h�,U�W���W�	K���1�\8�����-��1�l�c?�_mz5!Y�����B��_�7�}1�R��?󒜉��ٿʔ�jCl�':���*:��ФK�CU�Q��$]�ݮ���F
_�xOWq��;��l�2*��E��оJ\��-"������Z��|3N���a�09���ura�m�\�M�
A�i��E⑝;:_��z�Իޛ\�︮x��#U�R@�)������Y�dǭg.ĕ����a6��n��X�6��iY���������C�ծ�=0��N/��w|l1�!s95��4�����e�P*:��F��΢�����"��/��O��!?�H�.��0ž�Ia��ɲ�|�m0IgB�����}b�^,�)S_�j9�#��(E蟗)��\���@u[�����Ax��F�(�y�5��V���<�|��!��6t5ؔ�֏Ie�>�ڊ�{��t�0={���KBd�ݙ�[LVL�Dw��d��[K���(������_��H��ҷ�.c� ������3���( Vɉˋ��K���>v� Ӷ�>p�Ƞ�������բUm�&��o\�� }���*��Ώ:m�pĘ~���K �Zl�
�A`ZF (��l�j�������0#�.��t"%۞�L�|!
�C�e���@n����V����G;�L.룭M»��F�"�8&��8
�]:[�]sqc�8*�>�:������K+�R5
j��=��� �!��H|-,1o!��(��V�7����|�oo���m��*/a�'���	<����7c�>A\��s���3��ɏ|�.&߷�)��;�n?�w�k�o��
v���Y�&m.��i�&G����+=�V�8!��'%�p�ج�U��x��MQ�V:& ��H�	l��Ah�&��	�����TL��V����B�����1z�r��'��M�^��?g����y27�m�%/D� }�]3C�m{[o��095Xk�`cBC���O�!�w�Y�i*�3E�_m!�P��ƍ��^ �S�`��ߴ�h�}v���96?��	����wnTԟ	,�VL�W��"hL;�������7�Fg��SA1�U�$V�1$`,���E0.���> C��i��E��`�Gyѝ�B�O�}[A�哎��7Q�>�A�Ӓ �%u�|���q(��"�j>{�'��$w�^���W[�g!4��IE����l�*	��2�׶��Z�M�C�;:Ԁ��!°�-q���?>�h�Qf�slB��5f�o����$d>����`M��|ᙡ~����e%���*n%��VgW�J{"���[�5��7<hP�J��t��p_Dߏr�ݐ���=+��Dي� %���l����� �3���&�J�>$.��f��K	������#�ܮEu?��u��-�G!�7�"�L��qY(iC�z����}TCMa� �j���us����:�k��K 6o��K��N�p��%�,st|vW�FQ�����r{�^8;���+^����.|��U#zE5���g3��d+�����rZ��S7�Lc�Q�N#�o��0�:Cݬ?�4(k�'�Ll�3�������
˹ǒ��*dĒ)��_da����]����BS����>�'䩨)�y��j�⛿�}�U�
)_Kѧ�ʰ���L��!�;w���^)��w��K2>;�X�����/'�]wW�����J��诪�Hͅ��/�&�W�xl4T{B�ьίLx���{��92^Ф��.�@�������]�n�?�H�	��^�9���+��>d[���d�$�|��\u�@���]%��mA��ι|`��e/��S��+Ì�=�W��	�}|����e�#T2����{�[LbIT�|�Yf �c� ���I�����d�ܛ����X���X�8�4h�-�׶Y
�.,���'�Y�p�UZq%5�c�� ��ɶ��x��6�0���)Hɒ̉�gpgo7���a�8�!� �mx(��ROZXF�l�*5�#��Y��h���o ��Ե��Si7�(�ˤ���{����Z�����_��v�"�~,�y��Q{����A0Y���&o%�s��]]k/kU�^��B�ǀ5�̀C�f��LVS>�r�t$��uD^��Na��[��C��n{��vȡ�wf�8����},p�oe�:ƨ����X֝�ȨQ�=y
���{o�&D�N�+;l�(�Z'��ORq���X��	��͖��9�e�v�AOK
c�˕#�l���r��|3|�$��.��_tUs�=�Ԩ(J�yȻY�w��r{�u�8��
Pz�{4�� �ZG�1���g3��)�u	�������O/�@�W�%Λ��&g�#�U��g�7V
(��	�zP�S�z\ǋ ��y~����n�O�t�MĻ���ט[ٶvZq�OL��e�7/Z���Ε���V��}D8�s��wݮ`C.��n�CD;+^�?�>o	0�&��#7d����w��t��CҠ߲
�ƃ�u�h��`�OCM\�P֚+"B9��!��`:���U<|0���l��}�Od�sT�8	��:�}U���ȇ��)1v��p2_�ʗ{�&=gc!c͋�X,-���?����EN-l�b��x�!�4߅�F3`,Ҙq���%V�(�Bn�M}��-�&� ܲ%����;���4�%R,H-dٕx�|˽��{k���k����X�,C��8A������,�a�?�%���G���jҮi�S2)P��=�3P>���\�5�q��'!����m����+�dio�`C����-�1��Y�o�v��خ�}e�����g��~��7�h�|�{8�����mg��e�����1�B	�#�<��{,�/�6 ,(9�T7��ᣨt������c�*I|촪6�n��sQ��~ě$�>g5�s`n#~�����*���J,�eĿ=������Na�ʨ.�����Cy�:��u�����g��.?'o�|�t$΀�����D�fJ�4("kak2�MW����2��4�Y�U��m�8!�iK�c7#���l�3%�gD
JY�'�'=Ѣ!��(@$m��ڀS%�0t/�w�?)9��{��1-w�0[_��[·^��L�VG�I��D#�%qť�1����@rӗt����֨�#OՋD;IW�@��S�V,��y�5s��N�S�p-����wq��J����&'��8����[d{�8�r�G4;�3,�]A�o�^���� �	Xύ����D��Y�2!�l;��i��CN�X�7s��48͆J�����+��'�Ơ���o ��$P^d��$䆙Ϫ6f�s���S"˲QIq�b�]ȿEF��H����R;�+cޘ�d��o���OG����B�_�5��(>�.�X�^&���K�wD�;��a.�N\�6���sBcdj��O��ƚmލ�ݱ۠c��qߚp����ꮠ5�`_�	�1�l�j�(�}��۫V3�釁�Q����q�,�%�vԀ�| �Ю��_@]+��<V�c�eQxtɢ�N1+�)��I���a؝��S�&����j�7&ˬ��>|���%Z���K�ƍ��f�k|�F�/©�Y�ñ�ɴ�P��s��u���P^���穏|�'"jf_ZCf_2*��,w,���^���t
G������U�&!�iK��]&�I���_�`<��s
Q+	�o4�=����S��jv�1�P���BR�r9�������4ʍR�m��h!���A׊e�է�a�i� 9c�G�r)�?���Aa���%ϏPo�z�L�{��:��#M�(E�f�7qOU��'d���&��\�،(�)uױ5�����N�xؠ	+�� Y_�\�	���,_�b^�`�_��f����c^��o�""�彩OI����� Un�{.��Ǔ�s��P�l�2D��[�}mq=�r���I�v	�3�kJ�pM˛�����QN�.=ny�Q>�����0�3@�տ���L}
���o9�f}m��e�9�1G����_�|H�)����3"ec�q4�{!�����]�z�u��C�%��*�}�\�p�W�����!+F˶��.��Y57J��p�q��-벜�đ��>�7sd�t�k�K���gPd3�kVv8O��3ܪ�_D%������{�F� ߖ����Z�6�#��D��Gad�r~ti����p����b�<���u�_mErd�%�p|٫�L߲��
��X���m�τ�}�,ꁨ�gK�3e��J(\#\�>����i�E��=�%�v��rh�/(�+;�SW<*t�6O܏4ٚ:�KAu:�xV2�l4����'4:��+����
]�8S�OF����|�l^�&55L�3���	3e�Vuq\���&`<��\�7�AMɎg�	f�n+�+o9vc�9�3Qy�*-�J�*�+ˡ4�_��i�*�S���% ��%
�C)�J��r�}!)$�T1� e������s����g�����]�?��o�vA/�wg]/�,�c����
�]�w	A����K���Ұ�0Y���$f	�{�f؆+��Z'�����ҟ��Q�Z���4��=G��������8{�fxQ�hB3r������ z̸5��^����}
T�r�W�:�Y���r�2��曵-l�3�\���c�5W@�y���iY�K��Ua�d;N^����E�Ib�.=�rkjc���.��Ǘ���=!L^��'�4��0Ndp'�c]T�霄pj��:a.��`X΅M��*1��in�ϸ�~��i���GIO���ζ�}��3;�����>��!{�?�Ԣ࿢=r �Tk*�9�0�VڨJ�|�H[*�̬}���������A�C�,�	IR��/֌�4���W�iB����W� W`{	
�zB���&+sfxw���.	s_M��Q)��t������{�tQ���;�C�9����F�
 g.�D���H�T��!dB��J�.�v׾3͆Bk��=�3�����W8���|�᫗W,�N�H�q���|�U-}P�68e���n�5���x�V�A~�tj5!��F�r
g2:�?�Np�}�M��Bg� �r��9�0`0U�?�xv9*�n!���[�&f����\,�����k��.sYќW߈y�T}cG T�����;#�k�.��z�V����i�V67%�z8���mߍ�L�eQOU2|,�<��$�S����c�htl*�6�6���Рs3($ؽZ{�$v	�je��
nO!�5��T��*/(��X߂���]��Bt-�L|�\�$�<>����B ZF/��^�����&��T +@7/�����"h�R�@�,�$:J΁:b����M����
9(>6�;�F�,��6��`�_�C��_�_9/au�2�<M@w�XRM]\'B?d/4Q����J�j��7�e�r*�g�t\�^� z}�|�y��1#��*R�zMB_4�݂�D������R�%i����z}���&�D�6�2pd��`L>~4c�)Trc�[<MB�:A�����r=S}�<>�¶<E{�Ȫ\�K=��݂�]�x^�R�Db\B�̮�0Ү\�]�1q�YWq��T�HY�K[�)kcj�co���	}�!w��X�,dN"��}�{���k�#k�b�ؒ�a3��sX�S#��_6谿6eB3|���KfS��Y.�6��
	���]�+�Y�M �3�`p��o��R2��'�D!G�^�aF�� .W@�g�,2E�A�U�3q	iFo���(� �-�7�(: y���r���d����5�K�'wn*���z2�N䑑=ڷE+�p�ak��9���q�)���(�cBr2l�*��T���Ȇ�ۥɕ�mTuU`��H�l�..')���T�Ya>_/����'�ٟ�{���q�A�t�?L��!б�n����y���B�[�r䆵BȄ,dF�~Z�Y�E�\�$mc�%2'èR�S�
l�_��Y��`�!�rЗd����vˁ��L�c�9�o��]6;;g4����
z"M��P�R���2�ݦg^\k<����X[�����Ka������R��͠j5ܣ�#G�<k`�����$�!ˤ
țc]�]���룢𔚳�y�$ᎇ�b>�9�̳k�M(���]*�/B_8M?���hr��@T�����	�G���sG��QL�Gm�۬��U�:�/�����hÙzud�� z���p%��;>���aVQq�Y����̊V/᳡�G.��*Ņ�FY���5(`m��o6:�j�����͡�dŜFp��b�;_�8x0u�Z��G��*-�'Rڢ����/�Ϙ���I�!�Y�Y�,t� j����W�S%H�+h�<,�hbT�h����H�\Z�kO�0Q8��������?K5��54�]팻}@��c��f;@�k���hB��Du	��&��7<�T�l	��6P���
�3���6�'uU���*�M�*$�o�G�p.훃�2U��LoU'k`;�Y�h���ˬ�?e�8�Z����@���EẆ'�-��T���RA�3�F�YB�I�{(
41��"e��1���Xp�[^��t�����dd��\��1| �4p �I���� 7���v�Y�`uQX�Z+8$�.��M��,iz��x<*@H�Ϛ�S%�dX:F��L��P�q%x��T	�/���E��Q8�шI����8�;!���x@���y��g��:�%:V�-�𕑌�Y7Ϣ�ȷ�a9����5�j��L��N]Z?DLFܪ.��d������	^q��os/��mҢ��}�eT�}2�F��"�.�m��|:�af�Q�n>�hX��R:�E70�J��y )-$��ާk��C'
��.I5y����z�b�)�)/�*#�|����g��HF�|eҡ9l�#P�yc���dד��V��&qe
�ˮf��KT ��4�U�Zl?u%e���9rɁFi��G�H����rA��:���z�I�<�u���HfA�YGψ��_m�*�E��	��77�x�)�ens��T���O'������P�s����oy�y΂7�f6R�g��!����_*5辋җu-�ݐ�V�6M��h��Jׯ`�!� ��"�uw����[�
h�Qs}t���$�'�����q����~&B$4}�q��̷by�&2�yz*1�1��ą�M=t2�Cp�-Π��̤7á���f֦a�B�c�	&�.����X�2���Ax��ˢP�vO�%��e�!��jMs\'��K\���B�5�2��G��i�0�B�`ú�Q��nG�L�QA����MV�>�w�`��T��9��EX\2�!������'g���,��	0��t���i-�aO�;���f����t{|2K}ƷK�P14&��7W+��5Kc���`Cl!F�KW�S�ɵ�P�]�x�:ds��<�#��؄R^��Vz��Pż
�(|+����`�=߉�x�#}P��x��pd���I�Q񺪉�qe�����S�ß�U����@�v�*��&DDR��_�3F#�ͩ<�f5{���A��f�2�v=-�j7;��IT�{�A4�/�'�xv1z�}Vw��6'�jX7"��<IGPd~�ǯn=�0\��x�����h��6R�#\����8en��5��&k����$C{K^t��2^�+�����[$�4I��p��F"���r% �Zt���:/O�P�2��H�y�&q�}a"�0�+n�x{����L	`��
��˸z�2lζ�����w�$;ٓL���t��<_���~2W12/�־˼fߕw��H���KӋA�ڶ�p� ���C
�,�xC��������O�k`d�X����AZ�uh���iG@nZ1�2��!+:ix%%�;�F�θnE͗]y�]u��S�\>J9-1,�g���_b����c	({q})83�z#���kE/��T̂�f�n�]⭩�ˮ� ϡ$�ǋ����y!����+R��W�M��Q������Y���Q,/� ��y3)�g/�n���iŕ�L���/�/�V3��������I���猐6�_o.�	"^8�^ޢ�.}�s������§������;���_6��r�8��"�z��=��)U	5��kNzC���j����r��Ā��Sո�v�Y�a�)="�R�C�L[�yz͕��7N�>���\u6�v>{��F��6�G�`
8��-xq�Hy�	#}�"�ߠj4<�o\5̥�3?�����",f�h�mk��lab�	|�c椹�<fUM�(O~�g�l�G�:�B��D�/E����� &�l�//Ł ��r2���P ���`�}��4�xF�r�+㞚0��
�L��"�ۑL�c���B�o�G��qZ����8�OA��DRx�zwj
�=Tζ�(�ǽ�o%�ܧ�x�v�� hƒ�h㾪~�������O�Z@��r��� F��}��kC	�/c�UW��V��+�������[����.���3��/IK�[Zb����ߚw6G�2D��R�
{�m���Q`��k��b8H==OUW��V̮��~vS�������s��U¾*�/{�n� XkXܡ�dӚ�ʌ�u�܀�5c�wLuK��ŀ�J]eeFfW�6��l4Y�ޡϋv4 �I	s���`�GU�Xd�`�㌥�]����i��d;��VHF���"8r��q���3
\�'�Bʕ:'@�e��\K
� A���GcfKFV�6ȁ/�rLݾR�b��Ƭ�Să�{��X����y�Pk{`�J�]fp�����v�M�e���W����\�ٝ����6Ӓ7g�E�o�)�6����
�C4���q�8���ë���U�F����"�ߦJ̮S���T��r%���������r���т�l�;��r�u��玏��:ɝ�g%�7MI�uy�֛��9da�+9�wM���|�iV���`1H?��K��N3�����?8^�]��;@;ɽ@�M�(���J�R�\�X���� q� �J�R�Arhm�޵�U|rG	V+}�C$;��ڼ��
���Y����%gD*֣�%e����(�{�.,�ʽj$��;��,;c��I�%�ZO�=��N(�j�[���_2���h�W�1G�u�82�8N��(�1�$�״?����5��i��{$��� ]B�.��j���ˬ2F���͕�^Ha�������@h|�o{R��-�gӥ.��[`y�}�fGvf6�aٶZx�#	��*07J�E}o�p�q��ۉ�X-���4��SBM�(��Yc1�,���}j���R�v�p�ځ2|��\�=�������A����f}�^,�T�����6�3ǚ�U�/+ЩO��&tt�;�>U��x�}��v#|�����k*��ѡ�8([�M�?ǣ�1j��N>>�i.J
�@��*�&��fCĚsG0�-*Gu`��WF�R���l�hS�+��,3m����\���&_Ƥ�i�0εl[���
�2J��<cMJ��9c4�&5�k��ƻ�q�����6a)��|&bpoڷ2r�-}r�gpV�������{5z��u��T�v�a�[�;�z%��>�CV��M�k-aY��Q�H�F։�VII��3��2�c��w�t�)���W��wJ�-�s��o^?�WQ �B�/�
��6��~?)�~��jV� Z�	K��3���"�dK�>H���ێ�N�;
�C����7���;��F֤5W��-�P���q}�҄Iؓ�rWB�ث}�h�ИphX�}�=����`^
,�O�%f2�S��}��!��g�I���0���7
&�W��FO�v����?[Ѳ�~Sw�q1�,1�>HqB�e�ճ�W �/A��!�`���O���fV/~'b���T���C��hc�)%���"ex�Ln�����V	*����J\}Y��Z����<=Y��v��|���e������kBC_i�/q���E�,G�n�{ʷã�cka��+�	��b	.'F#��̡�NF=����s^4�Jԡyq����H�椩�ٓf��o OlAj�t�R�5����v�,uWt��MZ�%�}骍�̈�.Z���v�(;h����/����U���d|yDx��X3I?wY}�u��WN�"sL�u!�����F�β�ѡv�/�F���?-1���r9�΍3�_��c��@�`�(��baYHF��W��ΘH�HW~c�ԪVr")1�H��U_鷗l�qǟ��F�	표.��̛�k���0������,�c*t�#�o/&��+|Д��<��*+�1��}X隥'I��ף�#��D�~�K�*cRC1ɂ�X"�	6E��S�`�z�ޮ�U�n�н�b=���N�@�;>2�҈�A�����3/:_yF�����[���!Z��k�q(��;�-���+3����p:�z;�خT�
�+h{��[/Mܠ]iǁ_�X6�=�����S:�	���Q��#]��ҋf�%�� �@�x|U�ڼ��>$��'�i|���)`�^K �9>l����,����Vl��W>�ʁ�ļ������8�����?�K�*��"��A^�K/2��(X'/��5Y��Y��}-��F�tv����d�3�N�
̺L�z�ڮWcS�P�ö��J�D$�\�E��빾q�����Ja��O7�U����H����m�]b+k�=N֚]N�څj�N�����u�^���� E���J�/Qp!�M���JU°a�[�k�4�##d×l�+�����u?>���HJ�*_�[D�(*�a���贻��'j�������U�.3��K��%e)���[~��ޖO����:�#y��[�4N9�)t�Ԕ��"�PJک�9�<�.�UW���z�wA�%�T���՗wW�}&�W��ŵޭƣ�!��CU�
G���2���s�[w�J�;a��wDa��^�;�4U�r��������9F2����
 �`�������qt�gYJ�G����R��r5��#�������uԤ�OS,�犱�ey�>�/?�V�s���N��(�m���fpgᶐc��^�j�\S�Tl�d�l��M�I��1{j	4nL�mU2l#Q�Aa�H�1c�.�<o�@Z��&���o��S��E7���4��OS�=����v�����WO	9*�i��u[���j�tP�4���?�kʀ$����A�tڹ�r���+�+�1�s� K�ދ'�J��U�A�� V��H���t�0�\i��s�a���b��:�/Q�	��I��L���gap̈́&��_�Q��T�zY���+�"3��S9��۲!���h<� ��_����n���f�Y�������
��͉T#iy{��G��Vj%�ŗ��v'Z�q���X�-�Ʃrb��{�p�=�=.AF� �aQ�P���I;x�'���To����Bǋd}f�;�)�z �Sv�[ Z����l��M@�Y�H��pi�s�Ƴ��2�?şf�`�)M ���E�����d�~�
������m5��OcĬ$s��Π�6�	����~�^A(��x���p9�)-5_�1��3e�N��@GR:<�ե�[�$z�� Z��8�p�+�����w8mr��O��n��볕)��t��!,��*�OV�H�wG�xf��'s��ٯ�k�is�Ɵ�2Ti��|ʇb�>Tȯ�eXQ;�*Z��P�6��я���ſ�����e��X#�͢�u�,��l��,\�4N&�~��� �:ߜ��^��	�����<)r_��V��e�ϛ����8Y�E�$]���~.�wk7b���ȣ@F0eN�� �^�T2"��G$�c$T`�FSP��)��sFv_kR�����J����뫃 %�fH�~ϓ�.�� SNy���hm�����W�M���^��:@f�ۮ���_�J��l�"_ ���=z�T:��������۱B�P��i Q�D�WΧqL��L���h����9�a����w��LR�<�;x����A�y�*�Zלn$�S�E�.�#	5H	?��ߍTv�%y�nD��!��G��� �.�|�W��dB�T {�o�G�b#��-�(��ě��v͘�Q$�z�1Ux�;�e�VE�J���p���l����j[���U����"�ζ�[Q����G�ܶ�K�9"h0����9�¡���&eD�-���mV��8_��T��B��N��b[\u�Q�~%$�:����b��=��3���l���a��X�W&ϨV��D�c�1�>"�ZYk���Z�$5��?����=�~}�9
<o��g�l����6O��$r�nD�
�S��;%��z˄d��}��])r�u�'����YB�9����F!Ќ.�~��x:��S֮��_/.���>��b_4հ�Z�X�Û�<�v���1���A�9�.$��ի�}��e�1�u3*�֡���P.mq���O�\�fwki�k���g����
��%�u�i��������ڈ6��g�6�ة`	\����<Y�>) �nҎ��� ?Ѱ�p�%���塰�?�a�o��n�?�-T���* *���
-r�O|t��8�Rls�a�W�n��\!+�zg}��"L���?JOr�T�zߩd�X���s��x<~��<5�*���f����*����V�w(	
v%gq�^�){9���>E�ٮ���[6i�o�7Z- 9Z��1	�I��z@'b¤�-��"{���@����µ©��	UcA��}�d��ֲ�Ԯ��m��I��.Y��̓Q����p�Q``��rl&���O=8D�E���R�1\I8��m��^���#h���E���^����d1�<^�����������ȕ���t�4ځ��H���<�[��{����G�l���q_Nݟ�0�d�^�%���R�=�π���8��BI���u���\�%��K��K"P��@\�YI
�W�&mt��X����'>�X7�p�wP7nT��-��Q���4��ⵒ��Y�������M�SYji�o�1�.�>"3��x�`7$�~N�X������:��<S�GR����U<+�tV�PB�dF�8�m��񙩹;�Dq����2Z��b�����V�܈�cO��4;#u�Z��Q����M��wq���`9>�Ɲ��=�v6uuo$g���ݼe�A�!]c�s�c��M����	=6������EݛV�?��~��\�K&7�`O�0����6{OL��+~s^�XQ)9�/'Ʌa��V���">*f�/��>ֺd63]*��Po�l�vڕ��)g�o��Xf��ި�3sF��Î�r��U�A*F��ԇ���-zu�Z������I��#؎�7�`��q@Ή76|,HW���	��[�+��W�y���͋�Z�_�B�>Gq�p�C<���nQ�##����E���U���c�KJ���]_WF����q[v�6q�O@��YLa�/���;v[� �
lR[��>����Y��7��Z����O��/O�PΈU�",58�k��vQ�]��F���͜4r�"G��'�0�P�,�OY���F���q��H�; [�2��~]�P@α�&�f�����8�d5g�r_��ԁO�	��vZ(5�尻�f`e0���c_�,Oj��64�m��� '�����>����6�P� �l�.���̮Q+�I���:D�-����H��#��P@��8��A�;���"�8z-u��<p�rO�e�������wQ��q�)u|Al�+��Ӂ1VT�3,�	�0�W��T�![C3IWbV�f>��&��Wti9~B>M��c$�_e	u���2�Ez�T2�o ����ݹv���jn.���a�9���0�E^4egY?��*m��<z�}��Ч��tt��&�zt����wˁ��'�jV��l_nP£e�A}	�~����D#`��׈���l�)!�B��b��0<���n"�,񭿏�
���bH2��EM��$>���pj��@;�*�&g�H$�b�V���Eb��e-���[�Ȭ	v/)�ѫ|���{/��4HK����R���Q��5��~��k��������@��~Cts槡�g�N^/�����ڠ�s��'� ��B��P\�ܷ[��f�z�g��sy�َ��[��i�������QA#�6=�3�}����Y�E�Q�Z��!�1�t�Y��w��y:��/k]4�.��Xo@PdS�9܉`�'�'� ��x^$���\"M)i��RR}5_R�-X�F�1@&fQ]���EIш?��/]���!��)�����G=s�'̔��E�����*˄
�p�]�"o�ߛ��XK{U5��s�v.Y��0�����(s���^���&:�8>�ݦTj��%����VK�Eȑ�6��;��{^�몠Cyc�,.�f;��4��ٷ�j����~�Sj����xCvUD	��.3@��6D�ʰ%���'�p�M9����?&
�ss�P�z�zzhqO���*w�k���[���� }3yVj՜S�ԟEΛ ]a����N}�f��`?	�9��!�׀bu]��M*1G�ۦ�t-�������J�Gs_�J���e[��Ս�	�$Q�Q�y��s4�d_�%k��-`c�(P���������0G��ߧj�2UL�f�֤j)J���<�s���hd���w���:glk�Ge�.hV!��`=��T�H��ԯ�G0`���E4����\�X+� ���^�����AE��#fNN6<<�����#ݶ@�w�������.��9���ξ�5|��5r��}�j�q��CB�(3������ )w��GԒ
�@��`>�BM�Ư�d�s=����C�0)��d[��A2g�15�j��"֢�C���%?�9�iX �7S�B',�3-��茉��(���Ϭ��x�B�<LQ�U
%�M�4����6��ónrӫP�(h��AE�"�<ϲKa��{.d��0���\��Yf�i�i��⺭�zr�iI=��s���v����{��^r��D%�Ős�ψ�E�N]��/)c�kԿ؅/��r[6c�+J�n=�OQ�9ea]g���V"Y�LW6��a�%*0���o_���0����M����n�;��vB���1;of�,D�6�����5��+׳�1/�J4��J��fx5ô�UJ_>�0�����Z�����B�d��U[�>ѫ�����c;v�A�]2ݿ7�LBf�5Ʀ6�z�������:8T�뫜e�Zz�<�`��^�6'�Ng`�����y��xB���d׳8k�P
�/��ĸ����O�vH�] ���Ggi�U�/Z��FX��6H��~^�N��Xk��b��F�T�Eۿݾ������bs�ɺ/WO��}�-�^�W�u��r����%z��cD�mYR6��	�7�d���M��œ������%�R����ʹ� ᷱ@��O݇W��QU�ӎ�X�"�|+��V�NT
�S �c*��H��f ���Zc
yߢu������p�EJ���T)���Z�d�\��K�f��y�z��k�r��7���tv���Ax�H�_����p��X���	b�5����C��%� E�H
?)��!��lYG{�b���e�ɀ�e�I�Y~��O��m�q�3�R�=�M�njy:Nl�7��*����ƫ���(yS�����%��/�ja��d��MěxcGӮ≠$���1�̬o���ݞa9{��ۨ̀^T��u��;�� �y�b9��@>2�����將��~�8�t�Da�fO����奍�$�j�_��G�a�S��a���E����f� h��i��2)�h
��檁�����2�U6
��E��4��q��ٖ��G�T���;ڙ�%����89PxaS�+��U��ަ;�,5��چH��@�k�ꭁ��)��)aX����f$�|���)]�YA[g���^�1TK���Ň���"�R�r[6�gL�S��X@��y;���sH�#����r����8�q(�ɵb���H�(��͊+�e%l%�EaC�Pny�м�t�i�uݎfJ3�5r���5��(��_ݱ�K.� ��7��P�Y�t%��AM�`3{Z��1����X� ̦�fLWf)p�u��MsE:|���l�G<�44nR�����M�69Y��D��~uC�0ѻ5�r�n�y�
k�7� Q�n�MJ3�Ho���됉� 3�/��v� gO�Z�~��ɯ�6k�8rН�B��8�����*fP�����H̭�R󣮆J�܃'���o�d΃��b������G�?d�#t��Q߾�oU40�&\(qL�)9Nx�M�$�����["%�k�T��33 �Ȼ�c��9_;�����Û�&��hHJ�g�wj��Č|�6�.r��Fh#CZ��	����s�_~N�e:u{�9<�F?�Q(��W�+�Nu���!�?AV�Rm쇕O�B[�l�e������~w�����^H"{hq�~5H����0JO���/PE�xIfn
-<iH��y:���5�4�(���,���w� �p�7�����u�{EA����2����A� �h�y�?��%d�D@���C�^�s��!1:N�H5.�K3�-���0�Tbdb�,c{z�e�1�j����ڥ՟m2C�^Hr�K| ��]ݱ�ې��nv��tl�F��4����+.T�0�i����nE���;����?�L�MZQ�zz���~�x��h/82ë0f����:M�%���!?��ײ�D��Y�;���ξ_Ԍ4,^�OJ��Vg��0>dF�Y'
�DWj�X�Z�������"Z�f��[�k
��s�h�@��Jc�C�]�(g���r� �]Oզ^��:���HL��~��R�S:�سPg �ڧ-��(����]�s���N&�|;T�Ć�W��,B_�`��x��l"u+lϳ�L���C�e�簄x5�H�n�4Y����?#ެ6)<�W�[ˡ�}��Ű�x
��f:i����_�HT$x|���\~��$�l���5I��8��"paq����ٟd���8��2���n��+�a�&8N�*���}�>�dZ��V�/�X�m�w�N���j�y��ԠgoJB ����J!:V���eaŉ��A�W_����vh�	�rx@o��Tu�zؿ=�nS#��Mj�9E��U�PI�����;���&ֆ^ө�#Q�_~ 5Ad@�!2m��`���w�J9ᨏ2���<����mE7-$��"}e����^2��!�N3����U�����L<@�g�qj?�v���{u�q��*�����ZH'Kd��E�V3��{�,�!G��EV�n���p$V�?�"��Z���౉��Ӄ��mR��Oi�W��?�~օ��v���e�&�Xt����R��6��<#'3`j�{��X�h�*,]�W��5/���j�,�c��򝹘H�G�.(�x��k��1$0<H�@�r���L��@�����_���cu.�V �7���Θ"�.x]X6h$��|��R������
�5Cj{�m't�?]g-�����6#��]�@�}T/���pM[PzUݭgF<���F�@I��� e98�:iY��:�X���U����:3�`!����m��HE��W:�Q��Tyd"�'���9�5uĨÙ���lΰJ���45�m���!م\���8~��h41bp^_@�ڹ/^��]ޱ�(M?(�T*\l�h���/��~Nru5"?5�_D�[6����w���̕X!�EC����$�`��������/��a"p!������jǱ4ݚ!�0��.��("��� NtX�鲦�do&��\��ZBf�DD�<�����S��:�N{�&&1��7��4�g=1疥�쏭<� �a�(fOM־љ�\sg���N���KN�0�ܧ��2f�ۄ��&Uy�$���By�;r�$����t_��w�H�Qs����c���ϳ�e��p�G�8� ��z�/�Me�<������{�ry��FA�x}�*��	)u���K(Y?��l�C }'/Q�	Z�2s��|=�?��W+�9�t�0
`=$�K�O/��LF�&��I�Z�\1%�15����X��[ݪ�b53��a��d�J����YNٞ�Gq3!��^ͩ��a�]j~B��0h���SVVas��>-d���|��z���B%R���� H�ϬC%�m����@ �e�#H��T���m�2KFB ���g^[��x���F�=�A��t�g2��%��
�C��nL�@��M#����^��N/͎�˙���l����v-j\us�m�`�O��*[	��*o`�vQ&c�ح��)��?�!ȿ{?�Z�j��_t�H���cs�����˲D�\�߿�26�#��5�d�λs7���Ȇ9tΗՁ1�i�1��]C�G�Z
��f:f`��ʃ]��Mĭf�0��[mW���!�	P�I�{7�*]���8�0��7�F�ƀ�����*��-yE~5�يb��
�Y�ϖ����S�):l�� �/��K6:3}:��jo�V(�=��M��v�b�S	��*���覩3�<�~�V.��@��}���fGA���=#)��4s���r^�����7k޸���L�>џ���Y��3W}��������pf��'����vi�9&�L�#

�z�Q�[〉5v��7��B�{���\Z�vQ3i�ם�0�pOnHO0��A�N{�aDK�il5?������6_���IB����X�6�P9��}.�+f0y�����2+�:�Mc��l��kǙ�[��uaiz!��U!2���2�5l5��S������
9��o����q���@�$�8^9гTޯ��%��,s��_r�fi�slȐQ,3�kV��-U�q��	�����-�2�u��f�lAL��f2�u"��a6�2/%�/0�w������L{e��m]�3`��L��2�DHmd�6���"W[��oc�k{f�����l��r�=eT��9��^��b��Eb����{�������|��!9*��%Gs�I���is�����[_����:�����j-dS���]�rVB-��j�j�2��%ĩ��48# W�3;6}풑�#h���Ф�J�g1'l�ѪÔs%�z�����M��sŷ�/[5����b���)y���*� ?��~uK��d��	G3�ϝ/�&4����!�T��-��8O��ʨ>HC�okJ��D���p����1��f�KCn�vaYkă�`�Fh�~I5���={(���������4d&i�q��dɂ�4��,Dו�/����	��wޤ�Q�R���5���9���K���=w�1�-���H���A}�Y��s�������k�8�q��5�'�����U}t P!^5
>�._Yf-�35�G��Dq,�C\�^�Y��=�����itw끠8]P&��S8X��n�w�!v�P/��a�l�Ҷ�g��_�P���d�`+�la;\������+|��V���.�]�w
�[�Jڶ�Q�5�*���2@c���G�@�X�͎
b�!G�P����v���Bs����BY8��)y߱�ct8�����nr0y]}z0�6�S��$����I���U�hQ��������Vs�z�o㌫΁�cZ�ٺOM)��qI�<U�\���^������v��9� �͟3�������f���;FL�����S�!��{s<͓E����b�3���2�uuF�aCX�vxs��K��P:;F�C���w_'���n�(�s�,K̟��D5�ۜXK���+����JO�>������KQ��6�K��.P(Bj@�| �������șg��2{PY������_�+l>y?�1#K/6eF�,����>��s;��� �G��	��	2#��2i�+��4X��&�d@~R�1���_��d���j�V�����*���p�H�O�]�Al���00F@���冒bb�b�Q�(&8�֖	DH����_#ܬ���������0>����5hICśW�_O��C�}5�Sew�O��^[�s��ޡ;��r���mr�D����~0}�pʐ>:�8|�Y�no��5r�dU�T�C^�gF��E @�~��OJтJaxǰ����ߙ$�8�t�k�"}ma2�"=\~�~Ñ `����q ՝�0l�t��iH�i�$��g<.�����������2�/#k���`7띕u�n���3���kv?�p󱝤
��D�����V�$.S＝z���bU�-h�w@��i�����?�;`�%cb.싿�_V��T�M��q5ۙ`]ʃA�>��*Zy��U�̞>��H{^e}N�x2;�)5���-.�!�1�٢=S�a~	χ.n�4���9�ge�f'���EU< ����/M�_���c�06
�tN���y�xhv�1��ō�������r��B�-]@��d�r�Ƹ��=���Qɴ3���)�n�KNz�~t���6j��B���S.�y�w_��>ݯHu':e7,�*˚�dJzȵzcڰDy�tbi�`��A�e,�#qX�p�N�k
$��I�����k���K�]|��F*�7ፕ���d.t-8�����K�yXKB�&��{��B��UrЊ�����ӌJo�WQhA�^3�8��H+/N5+Ʈ8A�@�c�K�u����,���%�w������wܥ�;�ɳjڴ���l�%ϲ� q�` �4�~�m˂V�ꌙz�x���[��8y�3����WĖ
�H�H�hƭ�z;ox��T�����ٸte�y�$eo�:0�	�e����>��f���CE��ӂ�*,�M:́�r���
�5�3{G��Nư~Y5�6�r;������wkXY��K訢W���a]����ጄ�q̿<�|CjZ갃u�y?9����#~=�,��ҙ���k�� ���e�ٗ��.��= ��V��M�~o['��\�0��)#�(Q�_N�+2��w�־(`��h�_p��C~��g��K�����{�3V�y6�����h6�ez)��X�o�Ӈ���}T������1E�y�6�x�h�W����,7��*�+BJ}\�l��x�2`8*���0m	�I�>3I��b����Bg���
���3��P��x`M�v*�.*θO�������bV2�G�_��b}����}���9M���2���qB�Q��,C@!<@�_*�D\�������t?�f��6�8��F�U��D��I����a��_-H�9�xHCo̺m�;x�����#L�������GgYoA��IR�s��?���d�wx�0֞��a��8O�7�~��O��^���v=	l'����!��o�#�%��c�=]�P3n�����Z��!���!|��I��o���Wo�����ɤ��(���e���T�J��ڝ��Ə������LI���e��9��rs�6��B������^U.w\L���o|5�F�Q�(�[	b�s�Jck��,Rt���oG"�o���m�ǻNs�%����-SI�k�QU�c��M��ω)�1�$�M?���k8-ٱ�7�����4���S �9��L�����ݬ��р|�FN���LF_"������Q��6���r�Q8�	-͎Oi���Z�L�ӕ*Q��=���WU���wV7��r��d��8�?��V�R"y�ɰ����li�-�2���c	H��w�+7�|����b��F%�X~ �'`*���c�`�m[��!�P׹&�t���Q�Q	�Ng�[]���G��ҟ��S�#���6A���g7u��=�����@�V���
�d$��@�������7���u/�b�垩��XƨSi�kb^�pg,#����C�V3O�`O�@V�^ܿ���h��)�1
��hP?&_���U*F�u
�T>�oIY������E����Q����E _^f$��T>)zvip�",O2K^��j����'�39^-�FɦkL�&l��Z�Fp�SQNn���̣���1��� ��>y�A����a��3��^ڞ���Dچ�3�4�e�u�U�h7�tO?��؝񅖬2�z'�|�ʱh�Ew(�Rc*�|[�������
��� �D#po���"���}}4�t�u3� I�lҨ�9<��[����S�HP�F��a��q!xN\G�T��b~��w>4=.mګ��>��8�"��ˁ��R�<SH�E�B�L\�#�H�BT��^�~��2���Z]��"��eJ��~����!�	���w��sS�(�db���
�|��pL���^��>3sA� ���i����d��/u�vˡ�í0�N�7zu��#������w=��a����
x*�M�4����)��:-��Y�b�6\��0�n����MҲ�V�Ήj*�k��/o����h�d�t�H0�T%h�*�8�q�7��5���@{��wPo՜P�C���3��ZUix��5�Y	vp��:�O _q"F��v�a�w�܅}xE~��$�t�5�c�6m��/��c�P.ۙ�����IG�����"kR>��e	o$�!�H�Qy���KږC(�NP+�F���ڞ��k\�0�mpʋ
�>P׶1��AT��̹4���-A��'��|�q9��� �p	�Z���FR8��/�����h�mn!�ҙ
�F���v�;G;E��pu��: �r�^5-�zhX/� 'e_�s�ߩ� ՗�$�A���Qw���Nk���'ʒ��i<���@v/+NH����+S��R8aw)4U���H�ֽ��&�<��C�����!�VE>՟�]����͆C"��l�����*��ƥ��/j�Ctp';���9����ޣ�!c�3Y���&X�k��Mea���3�pt��;	��~}:�-�#Jy���T�\�ȓ�p��Z�T$��O�J����7JPP=If���l<Cv.�8��k��0?��0��@��^Jckp��h��\U���Dau4�_�tun�p^�z�Ձ�	ۓ���582@cm�č���bSd��iEHFv�C�s�W�XBz\
D�� ���Y\��ۺ�|�]SX�	�I�	��^���
�e�:�9�4�dB��z}xvr�1V��۞_�9E�̖�c֦o�	,��l��2�Z��2��wt1u�]�bʜW3�����<o�nj���*�AR�f������r�Q��7q�aQN_��M�my�A��Ojb��W�^9�F l^�_L�i�]�K�g�x��9qыI�Ĝ��8�]yL�o�KXuX�"��$A{�����)��e�q���`������j��8�I,��Xv���@d���2�Zoh��I��(�VP�	R[_(���m�iY�Hj�wK ����A��hk��]����M����VU]�|� �����;z���$<_����{I����~k�tf�*�y��t4�3��Y��q�B+9o�� ��8��yu�j��QR��G�_��[��\8�]w���V���X��{�3B_xX[Pe�:���
�&Ќ��S��l�Ƌ�BZm�Ɵڥ�R4��	��NyovǄ�+�P�U�����%I�� r7ߊ�|*�/(�)�f�
8q�#��U��aX̋�(�ʁt���L������&9o���]D-���� }��-�O��#���������E�[�]�+��_m�H��(�37PӘ�鐣�N7�s7�%V�\$�Ѣ��H�8��/�}&���~�<�?�g��,R�'>~�SN��j6��s��7�0$�����"����J� ����v�_8Q\�}#UA�����"P��;��|t%��8��v�+�!:i�(L�k��Z�u��07�����x�d�6w�܅���voOĶ9��)�_��.��r��ݩ��sΈ�1ef��7J"������}��d{��
��:�\����It�mybQEj����3=g�a�.���0�yq��˃v��^!a��j̨g�U܇�����%����ʍ�1"�<F��F7V��<�w:_c,L��x��Ϙ��L�&`�!\�qϜ���O���ړ�U4�5
���DZtt�$��[�>�GMt���Ԫ�:�'���0[���xYa���0�[7YkB�@�7
�4��N��ҙ��:�!�fg��Һ�7�h���L#��*ի� 8������Lj���?���V����"�]�Z��|��jRd��\�5�ro�C~��\��"v8�&�J�`�_\Qz��r�B'9�)O���I.�!�~0���G��m)HE�2���60�7��@{��Jt�ݡ��Ei���(�w��c��1�5f�[�xY���R�q�Խp4� �$�u�h?xq��[J*썩��n�J����8�� �׳��C�J���M������[&�c߳�uaZ�����C�W
�)7���p���S/h�ea����zb|Hܯz樂�Q��^��|[�$
�m
v�qk��ѝy�I}s���=�8�m7����-�6W k�=!����v�U�v�7?l#�?Q��3�ڰ�g���aU��z�f�u��G�:�(_J�K�H�RqS��� �����A�oJ���"J*������5�R$�K�灡bw?#��OiQF��+�V_͏IS1��-&˘o�{��.'��:L���q� -�Գ�3��\�ə�<�Ȳ��
�@^O���n�������{����,3��K��zX���Sဃ�p��%�۝Y�"`��U�d��S��^����B_��.:9�r�b,xNc��bY&9ćW#���!E���I6^|����H����ؽ�m���̭����>�Ob:�C�.I�*�v	s��}"g�X��Ohv��9µ6&C���-�W���>x�Bp'J�������Ӏ@���L�b�����ͨ��7�������q"/���\�������{��Mu%Q�rר��u�Y�~<�F�o:B�I3�h� #(��Ҙ�df�YBH�^I����SR�Ywm�Z��6m0CKD+濐9Lf����="`�����l�]#��a���)���/��TA"������2`�"�����Y��*����n��)��$����� :�}�ʀ	��{^����<V�p�n������4�z���CB����c&C�y�l䗿vʯ�3�l����G�8z0rWc�ؾ�����Nu5Y1��'ȸ@?I$��;)����^���=�s&$�;2ȣ�N���	�ͪ���cz�"tA�ĐF��,X���̹�_D�r����ˏ�����c"c`�&�`KDemԀ�N
�Z36�u�{����>���J���Ө���w�)e0�����wUn����L�G��r�'�.p�li�~�qEG�b
�J�e�Z֕�wH���r�����e19.dXr u9��h*�5��t�	oiS�bP��b)����=���L�����~�іg����Q~d�%G@M(�o�8(ݞ�Xfg2rA�~	
�t��zp1�.���R����|E,w����R ���ވ�H����o�H�t�d ~^O`�DG��0/'m������v��L�@��_>��m���U�+5������)��m��q��\�~Z���΍=�IA�Ȁ�kSf���.�1H0�;�X�;���3
���V?z�e��4tv�#� P&!�7	�>������оBnל����ebM�Kǉ��_�)��N� `�X��u���J���S3=>� k��$���0(N��5���gk��d����󛇲
RXc+��� ��@�	��Dd%f�Fd`������t{K���x� ���'���Dz���X[S$�8U�@��U;8�5��4��>���3���՘��v/bVj��,p.K�&�I��tp�lѠ��j��������AC¹Y)�a{�� �g�b���R�N�������e3]an����:N�����|�~��9��<���B��]��95�]j��ܦ��o�RqȲ���~b?��A�[�F}J�\�`3q%h�J�IQ��69�v�R�LL���?�pnH;�����k�	re�3�.����5օ1D�uٍ����&���6��H���UqP2zm�}�;j{���\� ��Bu�8�(�-��vV�UM�f$`�Y�WEZ�Zq�m�x+�گn�ǒ�!d��y�&DBt�Y1�K|�
Y�*`�?7�|5���!��l<�r�Q> ���̡�Du�����&�I]��7�O��M��!q&����(;��	!;������ �Z&�aN�X�$q#��!��ߎIs���\/����Q�@g�5U1쳅�q��(������=��n�o;���D�����sj(�/���j�����?��T a�����Wμ<�:E���m{/�Gʊ!�D���&d���6��r@�61)��"�;��+�`޴:��qU[[3������uNN���#��V��)��[�wZD�.�ٚ���e�۽�8z�>��f�h%#e�û�$��lw�I�R8.�c.՜V�x>����2�nO^um�3 �ec�:�>+�;׻�Z;r�jcuC��B�.u�WJޏ�E�|����e� ]v�V8>1����0���}�Ө��[�Kr[t?����w����0�h���2^<|�'�NaN����PO��Wq���z�����e�A_���3������b�2�n,�yP��f�_E��U𞡵���T/�/ڰS�o���ګ�5�}(nZ��K�kzJЛev���O��2��P�����KQwF�Z]Eŀ�Y
J�[w1�`g����c�C<�?r�&ٲd�"wU��
��������ץ�"�*6��xF�Hޣb� p-�/��r@�F�[�|��e�����O>�3��,���)Ul���$_}��OP�@����C愌�It�mO:�q��O�ǆ�V��B*D��Yħh���Ɂ�'���M�g�墯��z��=2���B��<�#�5d�#�F@*��NKP���y�$�{��6 /��u~ֲ�]��J*Y�4`�U8U��ZL@�Y�D\A���Ž�4P��< �
.�:�U�I�\N�M�:����R$,DnDHY��k�2`�e��͖�����������|��Ƞ��$�f�Y[�au�|��'H;�ڨ�4�roC�M�*�Q�s��� ���xv��w ������'i�	�ӊr��������L+!{�`����b��Qوo�蒳���5O�-�$��"�C��*QR�H:c9�lI4�=�w���De?�ȳ�0N ����1�(��qcyq���G3�Vۤ�T���ֈ5�ݼD�n'�)�UWh#�M��J-*3n]�~q2W*l�Swy�W��e]�8h'��8ۗ|9qz6�'���p_�g g�R����o@E~c7�������W*>��?�Չ�Wh\�i>��4P���Ϊ�oߏ鈧\�ů�R�M� ]�%��O����f*Ș�w�Ƹu ߝ�
�
�	a�Q�J����C�S�)����a:����)�ؤ���*Д�}�QOCu�>p3���ϡhb"d@�u�i��Jw���'� +�<
���ʵ��w��EMjd�In1J�&Ư�-����JMi}ʴ^d~Du��"�q�m]����hE� Ӻ������l�f�b�KH�Ll�@�� ���G-�o�.�bչk�4�M1-L
��˾M8�ґ>�J�q���Z�kL(�P�$)���?�$�G�
tL�L9�EF�24�����)�I�tz#YE��X�+�3�^�ѢJ(��;(�H�Az�D#qY`�{]��A���8+�v��|ɍ/y���S�Lt@oU���2�R�wY-L�`-�X�7}����H7��ȷ+Ka}e�q����v��gc�)��1�ޖ�[��jA���"<���͛D�xfJ����9|h�F��?=����k�nD�����I�J&`��<�@9?$inv�W���z�\Sw��'�g`��:�-ʠ-���PoO�7�k�j�ZH��3���?ʽ��u�#��}�T;A����2(3���&�����{�Y�k�����U[�#`c�P�Gl=�3�UB���-(:Ǣ�q��5�fmy��d���J�l8d�Q��6��R,��*� �N6�A]݀pPe�i�euj��'��u�"��`a�~bW�K��&#��$mr)/,s�
��L�NA����V-���eB����(uv����}�%������GPl�M����ȃ-�����[����=��.��u���ٶY���fg��,[��b�*6�����������*r[�\q��d=T_u�
������V�I�_��Ճ~8�>�^s��"ku���ST��P�����T+7��+u-�U0&�����ok�|�$�� Z��o){P���̙�	F5	-|sЋc�ȉz�
�"ոŶ��_�|�PY��x��מ�!s�1f��36�Pӹ8a �ԁɫ/'{����B-�?��ɏ�Ԟ���+�Lv0��r�"w4ZR�
	���XA�諾��W"�����C��V:n)	����(�^g��"[:ahqQ����Y5'g����M�G���QS��PXc�J�r�5�px(Jdu��f�~+����wEs��BK��ӥ���bg4�bH��0��� �[e�e{LeQ����p��v��/1�&�����@�H����'折�\g����t�<��)3�g��h'�eؤ��i����3{w̬��|��$Q2r�'��ч9]cbU��ؐu�)���}C3��w�6�e�O��
F��!w
"��ҙ��uM� u u�� ���a6�IO��g c�������j 3�����q�cY��:���l+	��&�_�;��7I(Y�=g�)�[HH�QAm�ٰ����Q�Դ�X�^#HR7a��s��9LXM�>s�k�H�-L?�X�|���dz�\?�p���f�➇�	*��*�??X�2������8��:��ƒ�R��*7Jv(I>j8mc��À�!wV���u7Q�̈́
>7%e���p�fS�����ٙ=��ĥ�]kh��Le�*�t�,2��Ou��_�t�j~�����ږީ��,w���2�L�M2���� �sƉ��B�s��Y�RC�o,l9��ԋ��v獠�ǹ�R�\_|�.�<�o9�qAC����L)(�4:$��y󒭫�����Z�t&���XSs�����sn�q�L<;�!dg��*8�<Y�ߣE�x�D_����J�ɳ��eTfb"o;!��ݸ��3w���h2$T�w��P��bS3�!u�_��{-�=CVf4+�fj0�����=���g"k3N>8�L���Qt���<�7�
�\g��?򴅉J���	�O�a�ġ�N�;,Gk������P�J�3���)�#2nn��L�:u������{����	ߨ���r���x�͆��;�0�	*���)Y�Hv�����PH~ݴ �x�
�u�D��u˒�N��Tfxy� �S�:��"�<gF[��CȦU��X��MO$����
O�g~EL�(e�����g~�#o=��y��7�?��z�rih�7��e��?(ڴ<D8��kP0 g5'����Yt�8n=�a�<p��@�e�+׫�s�w����|mw��=v)��.f���S�%My]�O����Y��PWփי�"̋H�{x��)��c��¬W�ʒV_�������͛���N.'� �e�Jr_ħgR�E�][]%vߏ̬�]g��^�� �T㡎{���M��;0o(��SJ�@��pF�0���u�/��k"��7*����8�;oƃ�L�>t��$(�3�Af �P���'`7T��i��X�X�2�x
# �r�������V0~�0��[�Ŕ�p(��oI�'�^@&p��������z TU�����-Ptb�Z}��]{��5;��!�e�s4�E�Gi8��SvU�_���,��%�u<v��6�)*_5�E�uȡXN$"��5����s��7.��a�tfW�*�3
ގ���UHY�7�RJ� ��#�}k���]��!��9�ߪ8���.]^(,���Z`�)|o����2쇲�'	��W���ΰ1���K���pU"~���-�"��M�"������mM>O�8��$IFJI��4u],a����8Ҙ��ZU/C]��M�����O7�l�QU��sL�2�RS�1 ��=f�����`����q��g�́!*!��&��*v$ƈ�1 qsFgBf��MIdwEU�� ��u�@�pD�0Z�3a��<�@Ty�^t s�;����vh��sÞW�f@���:H9�ʏ�u�0[�T�}5�`^4Z�ZG
)-�/w8��Ri#iH�H��ff�>��APЌ�C�[k3AݒNUUچ�+�#�(�#�b0_7��H�4��WX�|n��B%���T:S� 1�����tH��	S4�����w�|�U7���kk�F���5��
N�����o�q>�O�`g�� r"LT@) Yy�:����h�fHk4c<�<���)�r=k�fy9�9&Q|�B�g.�i��z��">�,[��A�,�ٹ�+哱�Wq���	�@Ma�x}��G���"�k%��7��c[�qL���~~��c�Âh@��-#T}ёpu##bls��Ϣ��I���6�}�V0�T��? �v�,��m.%��{8�3���5���o.��?&u��ʗ�^p�T�!Z�mb�(�1;Pd
�i���;�´߻�0����`��I~>�� ��hHqۚo�w�]>���3���DU-�$�(�4�szF4�T�?߯��jo`O(��A�n�\�QX�uH+Q]�5z_���KO
�|�,'Y�]2�ڢ�D�h�������;[�_ꖝT5׋�vk.��L���v�կ�?-PITR�N�3>kܚX�w?�P"Q��d�,����@�S\xU���H��{�P���d�������9��ꋸ��`�x���^ظ�u9�T՝���ׯEj������.c�T�a����4�I!�b���:�?��"���41�\�b%Ħ�I�H��� ����J.�+PN�*�㣔�z_�^�c�-((o�Z�/�(�ъ��b�^WmrIQQv�b��w����15ٜ��0�1���}^2z�fNC��r��d��t�I����v#�<�b)(p��.��U{`Ԉ�ɈR���(ƨW7���'uE�}���lA�)��@�n:#��(ܠC��v6��xԷ��v���bW��$c՜Y�������c-�X������mW��<<.TS��[o��2߆�ZU	�a�F�p�F��f���3=� ��g����nu���e�4qH�`��$8�Y�Ѥ���-���������_+��u���Պ���8t,��*��������}�/�2}���O���u���ؓ��R��Bo�8.�HW��R1��������4Z�q,���b�IG��O�P�����J��C0�-JlnD�]T��G����Ȣ�,/t	�&gHoWT�9�������j�̘Ը��8�Iy�&�Teh�<����1�I̺Ң�S��{��Q��[vb�޳טq��놞G�#ވ|�o�|�"��
UF`?p2�*�t���I�"���+��u���)w���ö2�C��,	L�b�X!����8E��\je����6�n�n��dT6ܞy=g�q�7,:�6˿<��8 �ڣ�����2k��~�֝hN8|\ /��W��n������lۊj��P�Mq�k΍c1�m?�с�����@�2��o���L^�����2x����σ�h���YG]ahH!(Dz��߳9"�S:�ָݜzg	�a��� �𓭄I����L�via�1z� ���P������3?�ߝ�.-�x�Ic�QZb����� �f[6v��^ %��_Sh��D�l����V����A��/)���,��ඩ&ibI
��W٬��l���[i����[�K	k�v�/���
��7>�yMxo��&F��~�](�Q����åػ��G�(�K�>t�x��t�=��H9fa=u�����'?�0�ϰ[/��w���۶(�W�:�<Z��o���=���P$`P�Ol�ѳ*�tW���&�p}�R��Vj�FUb��AH-֨d �:V��+��N5x���oIkQ�N����c�Qp�zc��i��Y��lư�mN�@��:���|MS�C(!
 ��f�,�z;9i5S+�����xI�t@����I��J,*,ՑA$S�,r��\��c�ع�u����7�V�W��?�VI�sW�ݬ5ŵ����26/[}1���V/��6�bd�1��HX�.�(����jYE�Q�(L���ffm���W���ڬR�i:��'�
j���+zm�ܕ��X�(Zr�ÅZ�0ڣ�B|�8KB�[����"b
n�w�o�Q#Q�ݣ��ϳ"��7S�j�C!g@��@W:xG\j@s(��=�mZ�_%/f��޵v����n�)�H�I���p9ؚ�8���2�b��'9�%mK�~�'H�����]��F������#��k�󢆂��l���_9̀�6V[} H@,$G��D����Q�o�Jۋ�D�!�'"�1Hإ���n
;���){�h�<��Ƭ��4U�o6�n��.Oܱ�7B����o�_;=?8�<*P�ϸ7Yl�p��ǐ���PSg��j��gm)�4F����4���9Q�=��`�c3�2'��Oi��T�vmr3�1�U"�v��B�=Q��ɱZ��TRi��-��q�)J@#�fhr�涁��j�Mu�x:����w�9������j&��K쓍f| aǽS�`-���wSڮt�ם��Z�2zdg�Yr�OA�\7-�$J��3b??�dU�����
�0V��� �UK���}�� Q��Xy?��M{���.R�h��(�� '�0;D#
��\�ʂa���>��ϝ�z��+���U^�.�*�3ĝ�������/�G����1��}*��	�Q���N���p��f9jpBO/�������<J8��|x%�R�-i�[޳`���;t$���c���l{G,�zQ %af���|�ZE�1��V~9����ׂ7�P 1�jI����9��gN�}_ ᤷ���=˓���l�64bћA����2��
��1AK�;&vo��$�:�iMm=R`����QASv��|�������حn�3E��W�U�ס;O�R>
��I 4���_�P�Y��MV)�쵶8���>��U9�m�Ti`����q
Ǿ'?G��"��h��F�P���{�9�T��TXK��e�f^�����{�^�ך
���:�Xڬ�